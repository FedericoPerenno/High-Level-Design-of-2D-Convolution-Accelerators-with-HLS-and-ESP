
//------> ./conv2dlb_cxx_catapult_ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> ./conv2dlb_cxx_catapult_ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> ./conv2dlb_cxx_catapult_ccs_sync_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2dlb_cxx_catapult_ccs_sync_out_wait_v1 (vld, irdy, ivld, rdy);
  parameter integer rscid = 1;

  input  ivld;
  output irdy;
  output vld;
  input  rdy;

  wire   irdy;
  wire   vld;

  assign vld = ivld;
  assign irdy = rdy;
endmodule

//------> /tools/calypto/CATAPULT_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./conv2dlb_cxx_catapult_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2dlb_cxx_catapult_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./conv2dlb_cxx_catapult_ccs_sync_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2dlb_cxx_catapult_ccs_sync_in_wait_v1 (rdy, vld, irdy, ivld);
  parameter integer rscid = 1;

  output rdy;
  input  vld;
  input  irdy;
  output ivld;

  wire   ivld;
  wire   rdy;

  assign ivld = vld;
  assign rdy = irdy;
endmodule

//------> ./conv2dlb_cxx_catapult_ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2dlb_cxx_catapult_ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0

    generate
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> ./conv2dlb_cxx_catapult_ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module esp_acc_conv2dlb_cxx_catapult_ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;  // clock enable polarity
    parameter integer ph_arst  = 1;  // async reset polarity
    parameter integer ph_srst  = 1;  // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd;
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
// synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      count = 32'b0;
      peak  = 32'b0;
    end
// synopsys translate_on
  wire din_rdy_drv  ;
  wire dout_vld_drv ;
    wire                 active;
    wire                 din_vld_int;
    wire                 hs_init;

    //assign din_rdy  = din_rdy_drv;    // dout_rdy | (~stat[0] & hs_init);   // original
    assign din_rdy = (fifo_sz > 0) ? (~stat[0] | dout_rdy) && hs_init : dout_rdy ;
    assign dout_vld = dout_vld_drv;
    assign is_idle = (~((din_vld && din_rdy) || (dout_vld && dout_rdy))) && hs_init;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
    assign din_vld_int = din_vld & hs_init;
    assign active =   (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);

      assign din_rdy_drv = dout_rdy | (~stat[0] & hs_init);
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign size_t = (count - {31'b0 , (dout_rdy & stat[fifo_sz-1])}) + { 31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use, no tx)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int  & (~dout_rdy)) // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          if (dout_rdy & stat_behind )
          begin
            // pop n shift
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_nxt & ~((~dout_rdy) & stat[i]))
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0))
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i)%8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]) | ~(active);
          end
        end

        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else
          count_t = n_elem[31:0];
        count = count_t;
// synopsys translate_off
        if ( peak < count )
          peak = count;
// synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      esp_acc_conv2dlb_cxx_catapult_ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        esp_acc_conv2dlb_cxx_catapult_ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        esp_acc_conv2dlb_cxx_catapult_ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
    end
    endgenerate

`ifdef RDY_ASRT
    generate
    if (ph_clk==1)
    begin: POS_CLK_ASSERT

       property rdyAsrt ;
         @(posedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Pos: assert property(rdyAsrt);

    end else if (ph_clk==0)
    begin: NEG_CLK_ASSERT

       property rdyAsrt ;
         @(negedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Neg: assert property(rdyAsrt);

    end
    endgenerate

`endif

endmodule



//------> ./conv2dlb_cxx_catapult_ccs_pipe_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 */

module esp_acc_conv2dlb_cxx_catapult_ccs_pipe_v5 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;

// synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = din_vld & !din_rdy;
    assign read_stall  = dout_rdy & !dout_vld;
// synopsys translate_on

    esp_acc_conv2dlb_cxx_catapult_ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld),
        .din_rdy  (din_rdy),
        .din      (din),
        .dout_vld (dout_vld),
        .dout_rdy (dout_rdy),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ./conv2dlb_cxx_catapult_ccs_sync_pipe_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2dlb_cxx_catapult_ccs_sync_pipe_v1 (dout_vld, dout_rdy, din_vld, din_rdy);
  parameter integer rscid = 1;

  input  din_vld;
  output dout_vld;
  input  dout_rdy;
  output din_rdy;

  wire   dout_vld;
  wire   din_rdy;

  assign dout_vld = din_vld;
  assign din_rdy = dout_rdy;
endmodule

//------> ./conv2dlb_cxx_catapult.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   perenno@esp
//  Generated date: Sat Nov 26 10:28:19 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_staller (
  clk, rst, core_wen, core_wten, config_done_cnsi_wen_comp, load_done_cnsi_wen_comp,
      compute_done_cnsi_wen_comp, store_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input config_done_cnsi_wen_comp;
  input load_done_cnsi_wen_comp;
  input compute_done_cnsi_wen_comp;
  input store_done_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = config_done_cnsi_wen_comp & load_done_cnsi_wen_comp & compute_done_cnsi_wen_comp
      & store_done_cnsi_wen_comp;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp
    (
  clk, rst, store_done_cnsi_oswt_unreg, store_done_cnsi_bawt, store_done_cnsi_wen_comp,
      store_done_cnsi_biwt, store_done_cnsi_bdwt, store_done_cnsi_bcwt
);
  input clk;
  input rst;
  input store_done_cnsi_oswt_unreg;
  output store_done_cnsi_bawt;
  output store_done_cnsi_wen_comp;
  input store_done_cnsi_biwt;
  input store_done_cnsi_bdwt;
  output store_done_cnsi_bcwt;
  reg store_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign store_done_cnsi_bawt = store_done_cnsi_biwt | store_done_cnsi_bcwt;
  assign store_done_cnsi_wen_comp = (~ store_done_cnsi_oswt_unreg) | store_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      store_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      store_done_cnsi_bcwt <= ~((~(store_done_cnsi_bcwt | store_done_cnsi_biwt))
          | store_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl
    (
  core_wen, store_done_cnsi_oswt_unreg, store_done_cnsi_iswt0, store_done_cnsi_ivld,
      store_done_cnsi_biwt, store_done_cnsi_bdwt, store_done_cnsi_bcwt, store_done_cnsi_irdy_core_sct
);
  input core_wen;
  input store_done_cnsi_oswt_unreg;
  input store_done_cnsi_iswt0;
  input store_done_cnsi_ivld;
  output store_done_cnsi_biwt;
  output store_done_cnsi_bdwt;
  input store_done_cnsi_bcwt;
  output store_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire store_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign store_done_cnsi_bdwt = store_done_cnsi_oswt_unreg & core_wen;
  assign store_done_cnsi_biwt = store_done_cnsi_ogwt & store_done_cnsi_ivld;
  assign store_done_cnsi_ogwt = store_done_cnsi_iswt0 & (~ store_done_cnsi_bcwt);
  assign store_done_cnsi_irdy_core_sct = store_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp
    (
  clk, rst, compute_done_cnsi_oswt_unreg, compute_done_cnsi_bawt, compute_done_cnsi_wen_comp,
      compute_done_cnsi_biwt, compute_done_cnsi_bdwt, compute_done_cnsi_bcwt
);
  input clk;
  input rst;
  input compute_done_cnsi_oswt_unreg;
  output compute_done_cnsi_bawt;
  output compute_done_cnsi_wen_comp;
  input compute_done_cnsi_biwt;
  input compute_done_cnsi_bdwt;
  output compute_done_cnsi_bcwt;
  reg compute_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign compute_done_cnsi_bawt = compute_done_cnsi_biwt | compute_done_cnsi_bcwt;
  assign compute_done_cnsi_wen_comp = (~ compute_done_cnsi_oswt_unreg) | compute_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      compute_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      compute_done_cnsi_bcwt <= ~((~(compute_done_cnsi_bcwt | compute_done_cnsi_biwt))
          | compute_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl
    (
  core_wen, compute_done_cnsi_oswt_unreg, compute_done_cnsi_iswt0, compute_done_cnsi_ivld,
      compute_done_cnsi_biwt, compute_done_cnsi_bdwt, compute_done_cnsi_bcwt, compute_done_cnsi_irdy_core_sct
);
  input core_wen;
  input compute_done_cnsi_oswt_unreg;
  input compute_done_cnsi_iswt0;
  input compute_done_cnsi_ivld;
  output compute_done_cnsi_biwt;
  output compute_done_cnsi_bdwt;
  input compute_done_cnsi_bcwt;
  output compute_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire compute_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign compute_done_cnsi_bdwt = compute_done_cnsi_oswt_unreg & core_wen;
  assign compute_done_cnsi_biwt = compute_done_cnsi_ogwt & compute_done_cnsi_ivld;
  assign compute_done_cnsi_ogwt = compute_done_cnsi_iswt0 & (~ compute_done_cnsi_bcwt);
  assign compute_done_cnsi_irdy_core_sct = compute_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp
    (
  clk, rst, load_done_cnsi_oswt_unreg, load_done_cnsi_bawt, load_done_cnsi_wen_comp,
      load_done_cnsi_biwt, load_done_cnsi_bdwt, load_done_cnsi_bcwt
);
  input clk;
  input rst;
  input load_done_cnsi_oswt_unreg;
  output load_done_cnsi_bawt;
  output load_done_cnsi_wen_comp;
  input load_done_cnsi_biwt;
  input load_done_cnsi_bdwt;
  output load_done_cnsi_bcwt;
  reg load_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign load_done_cnsi_bawt = load_done_cnsi_biwt | load_done_cnsi_bcwt;
  assign load_done_cnsi_wen_comp = (~ load_done_cnsi_oswt_unreg) | load_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      load_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      load_done_cnsi_bcwt <= ~((~(load_done_cnsi_bcwt | load_done_cnsi_biwt)) | load_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl
    (
  core_wen, load_done_cnsi_oswt_unreg, load_done_cnsi_iswt0, load_done_cnsi_irdy_core_psct,
      load_done_cnsi_ivld, load_done_cnsi_biwt, load_done_cnsi_bdwt, load_done_cnsi_bcwt,
      load_done_cnsi_irdy_core_sct
);
  input core_wen;
  input load_done_cnsi_oswt_unreg;
  input load_done_cnsi_iswt0;
  input load_done_cnsi_irdy_core_psct;
  input load_done_cnsi_ivld;
  output load_done_cnsi_biwt;
  output load_done_cnsi_bdwt;
  input load_done_cnsi_bcwt;
  output load_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire load_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign load_done_cnsi_bdwt = load_done_cnsi_oswt_unreg & core_wen;
  assign load_done_cnsi_biwt = load_done_cnsi_ogwt & load_done_cnsi_ivld;
  assign load_done_cnsi_ogwt = load_done_cnsi_iswt0 & (~ load_done_cnsi_bcwt);
  assign load_done_cnsi_irdy_core_sct = load_done_cnsi_irdy_core_psct & load_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp
    (
  clk, rst, config_done_cnsi_oswt_unreg, config_done_cnsi_bawt, config_done_cnsi_wen_comp,
      config_done_cnsi_biwt, config_done_cnsi_bdwt, config_done_cnsi_bcwt
);
  input clk;
  input rst;
  input config_done_cnsi_oswt_unreg;
  output config_done_cnsi_bawt;
  output config_done_cnsi_wen_comp;
  input config_done_cnsi_biwt;
  input config_done_cnsi_bdwt;
  output config_done_cnsi_bcwt;
  reg config_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign config_done_cnsi_bawt = config_done_cnsi_biwt | config_done_cnsi_bcwt;
  assign config_done_cnsi_wen_comp = (~ config_done_cnsi_oswt_unreg) | config_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      config_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      config_done_cnsi_bcwt <= ~((~(config_done_cnsi_bcwt | config_done_cnsi_biwt))
          | config_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl
    (
  core_wen, config_done_cnsi_oswt_unreg, config_done_cnsi_iswt0, config_done_cnsi_ivld,
      config_done_cnsi_biwt, config_done_cnsi_bdwt, config_done_cnsi_bcwt, config_done_cnsi_irdy_core_sct
);
  input core_wen;
  input config_done_cnsi_oswt_unreg;
  input config_done_cnsi_iswt0;
  input config_done_cnsi_ivld;
  output config_done_cnsi_biwt;
  output config_done_cnsi_bdwt;
  input config_done_cnsi_bcwt;
  output config_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire config_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign config_done_cnsi_bdwt = config_done_cnsi_oswt_unreg & core_wen;
  assign config_done_cnsi_biwt = config_done_cnsi_ogwt & config_done_cnsi_ivld;
  assign config_done_cnsi_ogwt = config_done_cnsi_iswt0 & (~ config_done_cnsi_bcwt);
  assign config_done_cnsi_irdy_core_sct = config_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp
    (
  clk, rst, acc_done_rsci_bawt, acc_done_rsci_biwt, acc_done_rsci_bdwt
);
  input clk;
  input rst;
  output acc_done_rsci_bawt;
  input acc_done_rsci_biwt;
  input acc_done_rsci_bdwt;


  // Interconnect Declarations
  reg acc_done_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign acc_done_rsci_bawt = acc_done_rsci_biwt | acc_done_rsci_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      acc_done_rsci_bcwt <= 1'b0;
    end
    else begin
      acc_done_rsci_bcwt <= ~((~(acc_done_rsci_bcwt | acc_done_rsci_biwt)) | acc_done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl
    (
  core_wen, acc_done_rsci_oswt_unreg, acc_done_rsci_iswt0, core_wten, acc_done_rsci_biwt,
      acc_done_rsci_bdwt
);
  input core_wen;
  input acc_done_rsci_oswt_unreg;
  input acc_done_rsci_iswt0;
  input core_wten;
  output acc_done_rsci_biwt;
  output acc_done_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign acc_done_rsci_bdwt = acc_done_rsci_oswt_unreg & core_wen;
  assign acc_done_rsci_biwt = (~ core_wten) & acc_done_rsci_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2dlb_cxx_catapult_config_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2dlb_cxx_catapult_config_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_staller (
  core_wen, conf_info_rsci_wen_comp, plm_conf_load_rsci_wen_comp, plm_conf_compute_rsci_wen_comp,
      plm_conf_store_rsci_wen_comp, done_rsci_wen_comp
);
  output core_wen;
  input conf_info_rsci_wen_comp;
  input plm_conf_load_rsci_wen_comp;
  input plm_conf_compute_rsci_wen_comp;
  input plm_conf_store_rsci_wen_comp;
  input done_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & plm_conf_load_rsci_wen_comp & plm_conf_compute_rsci_wen_comp
      & plm_conf_store_rsci_wen_comp & done_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt_unreg, done_rsci_bawt, done_rsci_wen_comp, done_rsci_biwt,
      done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bawt = done_rsci_biwt | done_rsci_bcwt;
  assign done_rsci_wen_comp = (~ done_rsci_oswt_unreg) | done_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt_unreg, done_rsci_iswt0, done_rsci_biwt, done_rsci_bdwt,
      done_rsci_bcwt, done_rsci_ivld_core_sct, done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt_unreg;
  input done_rsci_iswt0;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt_unreg & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_iswt0 & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_dp
    (
  clk, rst, plm_conf_store_rsci_oswt_unreg, plm_conf_store_rsci_bawt, plm_conf_store_rsci_wen_comp,
      plm_conf_store_rsci_biwt, plm_conf_store_rsci_bdwt, plm_conf_store_rsci_bcwt
);
  input clk;
  input rst;
  input plm_conf_store_rsci_oswt_unreg;
  output plm_conf_store_rsci_bawt;
  output plm_conf_store_rsci_wen_comp;
  input plm_conf_store_rsci_biwt;
  input plm_conf_store_rsci_bdwt;
  output plm_conf_store_rsci_bcwt;
  reg plm_conf_store_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_store_rsci_bawt = plm_conf_store_rsci_biwt | plm_conf_store_rsci_bcwt;
  assign plm_conf_store_rsci_wen_comp = (~ plm_conf_store_rsci_oswt_unreg) | plm_conf_store_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_store_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_conf_store_rsci_bcwt <= ~((~(plm_conf_store_rsci_bcwt | plm_conf_store_rsci_biwt))
          | plm_conf_store_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl
    (
  core_wen, plm_conf_store_rsci_oswt_unreg, plm_conf_store_rsci_iswt0, plm_conf_store_rsci_irdy,
      plm_conf_store_rsci_biwt, plm_conf_store_rsci_bdwt, plm_conf_store_rsci_bcwt,
      plm_conf_store_rsci_ivld_core_sct
);
  input core_wen;
  input plm_conf_store_rsci_oswt_unreg;
  input plm_conf_store_rsci_iswt0;
  input plm_conf_store_rsci_irdy;
  output plm_conf_store_rsci_biwt;
  output plm_conf_store_rsci_bdwt;
  input plm_conf_store_rsci_bcwt;
  output plm_conf_store_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire plm_conf_store_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_store_rsci_bdwt = plm_conf_store_rsci_oswt_unreg & core_wen;
  assign plm_conf_store_rsci_biwt = plm_conf_store_rsci_ogwt & plm_conf_store_rsci_irdy;
  assign plm_conf_store_rsci_ogwt = plm_conf_store_rsci_iswt0 & (~ plm_conf_store_rsci_bcwt);
  assign plm_conf_store_rsci_ivld_core_sct = plm_conf_store_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp
    (
  clk, rst, plm_conf_compute_rsci_oswt_unreg, plm_conf_compute_rsci_bawt, plm_conf_compute_rsci_wen_comp,
      plm_conf_compute_rsci_biwt, plm_conf_compute_rsci_bdwt, plm_conf_compute_rsci_bcwt
);
  input clk;
  input rst;
  input plm_conf_compute_rsci_oswt_unreg;
  output plm_conf_compute_rsci_bawt;
  output plm_conf_compute_rsci_wen_comp;
  input plm_conf_compute_rsci_biwt;
  input plm_conf_compute_rsci_bdwt;
  output plm_conf_compute_rsci_bcwt;
  reg plm_conf_compute_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_compute_rsci_bawt = plm_conf_compute_rsci_biwt | plm_conf_compute_rsci_bcwt;
  assign plm_conf_compute_rsci_wen_comp = (~ plm_conf_compute_rsci_oswt_unreg) |
      plm_conf_compute_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_compute_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_conf_compute_rsci_bcwt <= ~((~(plm_conf_compute_rsci_bcwt | plm_conf_compute_rsci_biwt))
          | plm_conf_compute_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl
    (
  core_wen, plm_conf_compute_rsci_oswt_unreg, plm_conf_compute_rsci_iswt0, plm_conf_compute_rsci_irdy,
      plm_conf_compute_rsci_biwt, plm_conf_compute_rsci_bdwt, plm_conf_compute_rsci_bcwt,
      plm_conf_compute_rsci_ivld_core_sct
);
  input core_wen;
  input plm_conf_compute_rsci_oswt_unreg;
  input plm_conf_compute_rsci_iswt0;
  input plm_conf_compute_rsci_irdy;
  output plm_conf_compute_rsci_biwt;
  output plm_conf_compute_rsci_bdwt;
  input plm_conf_compute_rsci_bcwt;
  output plm_conf_compute_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire plm_conf_compute_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_compute_rsci_bdwt = plm_conf_compute_rsci_oswt_unreg & core_wen;
  assign plm_conf_compute_rsci_biwt = plm_conf_compute_rsci_ogwt & plm_conf_compute_rsci_irdy;
  assign plm_conf_compute_rsci_ogwt = plm_conf_compute_rsci_iswt0 & (~ plm_conf_compute_rsci_bcwt);
  assign plm_conf_compute_rsci_ivld_core_sct = plm_conf_compute_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_dp
    (
  clk, rst, plm_conf_load_rsci_oswt_unreg, plm_conf_load_rsci_bawt, plm_conf_load_rsci_wen_comp,
      plm_conf_load_rsci_biwt, plm_conf_load_rsci_bdwt, plm_conf_load_rsci_bcwt
);
  input clk;
  input rst;
  input plm_conf_load_rsci_oswt_unreg;
  output plm_conf_load_rsci_bawt;
  output plm_conf_load_rsci_wen_comp;
  input plm_conf_load_rsci_biwt;
  input plm_conf_load_rsci_bdwt;
  output plm_conf_load_rsci_bcwt;
  reg plm_conf_load_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_load_rsci_bawt = plm_conf_load_rsci_biwt | plm_conf_load_rsci_bcwt;
  assign plm_conf_load_rsci_wen_comp = (~ plm_conf_load_rsci_oswt_unreg) | plm_conf_load_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_load_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_conf_load_rsci_bcwt <= ~((~(plm_conf_load_rsci_bcwt | plm_conf_load_rsci_biwt))
          | plm_conf_load_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl
    (
  core_wen, plm_conf_load_rsci_oswt_unreg, plm_conf_load_rsci_iswt0, plm_conf_load_rsci_irdy,
      plm_conf_load_rsci_biwt, plm_conf_load_rsci_bdwt, plm_conf_load_rsci_bcwt,
      plm_conf_load_rsci_ivld_core_sct
);
  input core_wen;
  input plm_conf_load_rsci_oswt_unreg;
  input plm_conf_load_rsci_iswt0;
  input plm_conf_load_rsci_irdy;
  output plm_conf_load_rsci_biwt;
  output plm_conf_load_rsci_bdwt;
  input plm_conf_load_rsci_bcwt;
  output plm_conf_load_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire plm_conf_load_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_load_rsci_bdwt = plm_conf_load_rsci_oswt_unreg & core_wen;
  assign plm_conf_load_rsci_biwt = plm_conf_load_rsci_ogwt & plm_conf_load_rsci_irdy;
  assign plm_conf_load_rsci_ogwt = plm_conf_load_rsci_iswt0 & (~ plm_conf_load_rsci_bcwt);
  assign plm_conf_load_rsci_ivld_core_sct = plm_conf_load_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_dp
    (
  clk, rst, conf_info_rsci_oswt_unreg, conf_info_rsci_bawt, conf_info_rsci_wen_comp,
      conf_info_rsci_idat_mxwt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  output conf_info_rsci_wen_comp;
  output [255:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  reg [255:0] conf_info_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bawt = conf_info_rsci_biwt | conf_info_rsci_bcwt;
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt_unreg) | conf_info_rsci_bawt;
  assign conf_info_rsci_idat_mxwt = MUX_v_256_2_2(conf_info_rsci_idat, conf_info_rsci_idat_bfwt,
      conf_info_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt <= conf_info_rsci_idat;
    end
  end

  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt_unreg, conf_info_rsci_iswt0, conf_info_rsci_biwt,
      conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt_unreg & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_iswt0 & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_12_14_32_10368_10368_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_12_14_32_10368_10368_32_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input clken_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_core_fsm (
  clk, rst, core_wen, fsm_output, LOAD_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input core_wen;
  output [3:0] fsm_output;
  reg [3:0] fsm_output;
  input LOAD_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_conv2dlb_cxx_catapult_load_core_core_fsm_1
  parameter
    core_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    LOAD_BATCH_LOOP_C_0 = 2'd2,
    main_C_1 = 2'd3;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2dlb_cxx_catapult_load_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 4'b0010;
        state_var_NS = LOAD_BATCH_LOOP_C_0;
      end
      LOAD_BATCH_LOOP_C_0 : begin
        fsm_output = 4'b0100;
        if ( LOAD_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = LOAD_BATCH_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 4'b1000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 4'b0001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_staller (
  clk, rst, core_wen, core_wten, conf_info_rsci_wen_comp, buf_linear_rsci_wen_comp,
      plm_kernel_rsci_wen_comp, dma_read_chnl_rsci_wen_comp, done_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input conf_info_rsci_wen_comp;
  input buf_linear_rsci_wen_comp;
  input plm_kernel_rsci_wen_comp;
  input dma_read_chnl_rsci_wen_comp;
  input done_rsci_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & buf_linear_rsci_wen_comp & plm_kernel_rsci_wen_comp
      & dma_read_chnl_rsci_wen_comp & done_rsci_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_dp
    (
  clk, rst, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2
);
  input clk;
  input rst;
  input [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt;
  output [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2;


  // Interconnect Declarations
  reg LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt;
  reg LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt_1;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt = LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt
      | LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt = MUX_v_32_2_2(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_bfwt, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt_1);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt <= 1'b0;
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt <= ~((~(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt
          | LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt)) | LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt);
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt_1 <= ~((~(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bcwt_1
          | LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1)) | LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1 ) begin
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_bfwt <= LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_ctrl
    (
  core_wen, core_wten, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_core_sct_pff, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_core_sct_pff;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt = LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg
      & core_wen;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt = (~ core_wten) & LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2 = LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1
      & core_wen;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1 = (~ core_wten) & LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_core_sct_pff = LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff
      & core_wen;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct
      = LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt, done_rsci_wen_comp, done_rsci_biwt, done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_wen_comp = (~ done_rsci_oswt) | done_rsci_biwt | done_rsci_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt, done_rsci_biwt, done_rsci_bdwt, done_rsci_bcwt, done_rsci_ivld_core_sct,
      done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_oswt & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
    (
  clk, rst, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_bawt, dma_read_chnl_rsci_wen_comp,
      dma_read_chnl_rsci_idat_mxwt, dma_read_chnl_rsci_biwt, dma_read_chnl_rsci_bdwt,
      dma_read_chnl_rsci_bcwt, dma_read_chnl_rsci_idat
);
  input clk;
  input rst;
  input dma_read_chnl_rsci_oswt_unreg;
  output dma_read_chnl_rsci_bawt;
  output dma_read_chnl_rsci_wen_comp;
  output [31:0] dma_read_chnl_rsci_idat_mxwt;
  input dma_read_chnl_rsci_biwt;
  input dma_read_chnl_rsci_bdwt;
  output dma_read_chnl_rsci_bcwt;
  reg dma_read_chnl_rsci_bcwt;
  input [63:0] dma_read_chnl_rsci_idat;


  // Interconnect Declarations
  reg [31:0] dma_read_chnl_rsci_idat_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_rsci_bawt = dma_read_chnl_rsci_biwt | dma_read_chnl_rsci_bcwt;
  assign dma_read_chnl_rsci_wen_comp = (~ dma_read_chnl_rsci_oswt_unreg) | dma_read_chnl_rsci_bawt;
  assign dma_read_chnl_rsci_idat_mxwt = MUX_v_32_2_2((dma_read_chnl_rsci_idat[31:0]),
      dma_read_chnl_rsci_idat_bfwt_31_0, dma_read_chnl_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_read_chnl_rsci_bcwt <= ~((~(dma_read_chnl_rsci_bcwt | dma_read_chnl_rsci_biwt))
          | dma_read_chnl_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_rsci_idat_bfwt_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( dma_read_chnl_rsci_biwt ) begin
      dma_read_chnl_rsci_idat_bfwt_31_0 <= dma_read_chnl_rsci_idat[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
    (
  core_wen, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_iswt0, dma_read_chnl_rsci_biwt,
      dma_read_chnl_rsci_bdwt, dma_read_chnl_rsci_bcwt, dma_read_chnl_rsci_irdy_core_sct,
      dma_read_chnl_rsci_ivld
);
  input core_wen;
  input dma_read_chnl_rsci_oswt_unreg;
  input dma_read_chnl_rsci_iswt0;
  output dma_read_chnl_rsci_biwt;
  output dma_read_chnl_rsci_bdwt;
  input dma_read_chnl_rsci_bcwt;
  output dma_read_chnl_rsci_irdy_core_sct;
  input dma_read_chnl_rsci_ivld;


  // Interconnect Declarations
  wire dma_read_chnl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_rsci_bdwt = dma_read_chnl_rsci_oswt_unreg & core_wen;
  assign dma_read_chnl_rsci_biwt = dma_read_chnl_rsci_ogwt & dma_read_chnl_rsci_ivld;
  assign dma_read_chnl_rsci_ogwt = dma_read_chnl_rsci_iswt0 & (~ dma_read_chnl_rsci_bcwt);
  assign dma_read_chnl_rsci_irdy_core_sct = dma_read_chnl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
    (
  clk, rst, dma_read_ctrl_rsci_bawt, dma_read_ctrl_rsci_irdy_mxwt, dma_read_ctrl_rsci_irdy,
      dma_read_ctrl_rsci_biwt, dma_read_ctrl_rsci_bdwt
);
  input clk;
  input rst;
  output dma_read_ctrl_rsci_bawt;
  output dma_read_ctrl_rsci_irdy_mxwt;
  input dma_read_ctrl_rsci_irdy;
  input dma_read_ctrl_rsci_biwt;
  input dma_read_ctrl_rsci_bdwt;


  // Interconnect Declarations
  reg dma_read_ctrl_rsci_bcwt;
  reg dma_read_ctrl_rsci_irdy_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_rsci_bawt = dma_read_ctrl_rsci_biwt | dma_read_ctrl_rsci_bcwt;
  assign dma_read_ctrl_rsci_irdy_mxwt = MUX_s_1_2_2(dma_read_ctrl_rsci_irdy, dma_read_ctrl_rsci_irdy_bfwt,
      dma_read_ctrl_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_rsci_bcwt <= ~((~(dma_read_ctrl_rsci_bcwt | dma_read_ctrl_rsci_biwt))
          | dma_read_ctrl_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_irdy_bfwt <= 1'b0;
    end
    else if ( dma_read_ctrl_rsci_biwt ) begin
      dma_read_ctrl_rsci_irdy_bfwt <= dma_read_ctrl_rsci_irdy;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
    (
  core_wen, core_wten, dma_read_ctrl_rsci_oswt_unreg, dma_read_ctrl_rsci_iswt0, dma_read_ctrl_rsci_biwt,
      dma_read_ctrl_rsci_bdwt
);
  input core_wen;
  input core_wten;
  input dma_read_ctrl_rsci_oswt_unreg;
  input dma_read_ctrl_rsci_iswt0;
  output dma_read_ctrl_rsci_biwt;
  output dma_read_ctrl_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_rsci_bdwt = dma_read_ctrl_rsci_oswt_unreg & core_wen;
  assign dma_read_ctrl_rsci_biwt = (~ core_wten) & dma_read_ctrl_rsci_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci_plm_kernel_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci_plm_kernel_wait_dp
    (
  clk, rst, plm_kernel_rsci_oswt_unreg, plm_kernel_rsci_bawt, plm_kernel_rsci_wen_comp,
      plm_kernel_rsci_biwt, plm_kernel_rsci_bdwt, plm_kernel_rsci_bcwt
);
  input clk;
  input rst;
  input plm_kernel_rsci_oswt_unreg;
  output plm_kernel_rsci_bawt;
  output plm_kernel_rsci_wen_comp;
  input plm_kernel_rsci_biwt;
  input plm_kernel_rsci_bdwt;
  output plm_kernel_rsci_bcwt;
  reg plm_kernel_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_kernel_rsci_bawt = plm_kernel_rsci_biwt | plm_kernel_rsci_bcwt;
  assign plm_kernel_rsci_wen_comp = (~ plm_kernel_rsci_oswt_unreg) | plm_kernel_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_kernel_rsci_bcwt <= ~((~(plm_kernel_rsci_bcwt | plm_kernel_rsci_biwt))
          | plm_kernel_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci_plm_kernel_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci_plm_kernel_wait_ctrl
    (
  core_wen, plm_kernel_rsci_oswt_unreg, plm_kernel_rsci_iswt0, plm_kernel_rsci_irdy,
      plm_kernel_rsci_biwt, plm_kernel_rsci_bdwt, plm_kernel_rsci_bcwt, plm_kernel_rsci_ivld_core_sct
);
  input core_wen;
  input plm_kernel_rsci_oswt_unreg;
  input plm_kernel_rsci_iswt0;
  input plm_kernel_rsci_irdy;
  output plm_kernel_rsci_biwt;
  output plm_kernel_rsci_bdwt;
  input plm_kernel_rsci_bcwt;
  output plm_kernel_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire plm_kernel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_kernel_rsci_bdwt = plm_kernel_rsci_oswt_unreg & core_wen;
  assign plm_kernel_rsci_biwt = plm_kernel_rsci_ogwt & plm_kernel_rsci_irdy;
  assign plm_kernel_rsci_ogwt = plm_kernel_rsci_iswt0 & (~ plm_kernel_rsci_bcwt);
  assign plm_kernel_rsci_ivld_core_sct = plm_kernel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci_buf_linear_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci_buf_linear_wait_dp
    (
  clk, rst, buf_linear_rsci_oswt_unreg, buf_linear_rsci_bawt, buf_linear_rsci_wen_comp,
      buf_linear_rsci_biwt, buf_linear_rsci_bdwt, buf_linear_rsci_bcwt
);
  input clk;
  input rst;
  input buf_linear_rsci_oswt_unreg;
  output buf_linear_rsci_bawt;
  output buf_linear_rsci_wen_comp;
  input buf_linear_rsci_biwt;
  input buf_linear_rsci_bdwt;
  output buf_linear_rsci_bcwt;
  reg buf_linear_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign buf_linear_rsci_bawt = buf_linear_rsci_biwt | buf_linear_rsci_bcwt;
  assign buf_linear_rsci_wen_comp = (~ buf_linear_rsci_oswt_unreg) | buf_linear_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_bcwt <= 1'b0;
    end
    else begin
      buf_linear_rsci_bcwt <= ~((~(buf_linear_rsci_bcwt | buf_linear_rsci_biwt))
          | buf_linear_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci_buf_linear_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci_buf_linear_wait_ctrl
    (
  core_wen, buf_linear_rsci_oswt_unreg, buf_linear_rsci_iswt0, buf_linear_rsci_irdy,
      buf_linear_rsci_biwt, buf_linear_rsci_bdwt, buf_linear_rsci_bcwt, buf_linear_rsci_ivld_core_sct
);
  input core_wen;
  input buf_linear_rsci_oswt_unreg;
  input buf_linear_rsci_iswt0;
  input buf_linear_rsci_irdy;
  output buf_linear_rsci_biwt;
  output buf_linear_rsci_bdwt;
  input buf_linear_rsci_bcwt;
  output buf_linear_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire buf_linear_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign buf_linear_rsci_bdwt = buf_linear_rsci_oswt_unreg & core_wen;
  assign buf_linear_rsci_biwt = buf_linear_rsci_ogwt & buf_linear_rsci_irdy;
  assign buf_linear_rsci_ogwt = buf_linear_rsci_iswt0 & (~ buf_linear_rsci_bcwt);
  assign buf_linear_rsci_ivld_core_sct = buf_linear_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_dp (
  clk, rst, conf_info_rsci_oswt, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt,
      conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt;
  output conf_info_rsci_wen_comp;
  output [231:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  reg [231:0] conf_info_rsci_idat_bfwt_231_0;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt) | conf_info_rsci_biwt
      | conf_info_rsci_bcwt;
  assign conf_info_rsci_idat_mxwt = MUX_v_232_2_2((conf_info_rsci_idat[231:0]), conf_info_rsci_idat_bfwt_231_0,
      conf_info_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt_231_0 <= conf_info_rsci_idat[231:0];
    end
  end

  function automatic [231:0] MUX_v_232_2_2;
    input [231:0] input_0;
    input [231:0] input_1;
    input [0:0] sel;
    reg [231:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_232_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_oswt & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_staller (
  core_wen, conf_info_rsci_wen_comp, buf_linear_rsci_wen_comp, plm_kernel_rsci_wen_comp,
      var_output_rsci_wen_comp, done_rsci_wen_comp
);
  output core_wen;
  input conf_info_rsci_wen_comp;
  input buf_linear_rsci_wen_comp;
  input plm_kernel_rsci_wen_comp;
  input var_output_rsci_wen_comp;
  input done_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & buf_linear_rsci_wen_comp & plm_kernel_rsci_wen_comp
      & var_output_rsci_wen_comp & done_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt_unreg, done_rsci_bawt, done_rsci_wen_comp, done_rsci_biwt,
      done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bawt = done_rsci_biwt | done_rsci_bcwt;
  assign done_rsci_wen_comp = (~ done_rsci_oswt_unreg) | done_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt_unreg, done_rsci_iswt0, done_rsci_biwt, done_rsci_bdwt,
      done_rsci_bcwt, done_rsci_ivld_core_sct, done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt_unreg;
  input done_rsci_iswt0;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt_unreg & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_iswt0 & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci_var_output_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci_var_output_wait_dp
    (
  clk, rst, var_output_rsci_oswt_unreg, var_output_rsci_bawt, var_output_rsci_wen_comp,
      var_output_rsci_biwt, var_output_rsci_bdwt, var_output_rsci_bcwt
);
  input clk;
  input rst;
  input var_output_rsci_oswt_unreg;
  output var_output_rsci_bawt;
  output var_output_rsci_wen_comp;
  input var_output_rsci_biwt;
  input var_output_rsci_bdwt;
  output var_output_rsci_bcwt;
  reg var_output_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign var_output_rsci_bawt = var_output_rsci_biwt | var_output_rsci_bcwt;
  assign var_output_rsci_wen_comp = (~ var_output_rsci_oswt_unreg) | var_output_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      var_output_rsci_bcwt <= 1'b0;
    end
    else begin
      var_output_rsci_bcwt <= ~((~(var_output_rsci_bcwt | var_output_rsci_biwt))
          | var_output_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci_var_output_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci_var_output_wait_ctrl
    (
  core_wen, var_output_rsci_oswt_unreg, var_output_rsci_iswt0, var_output_rsci_irdy,
      var_output_rsci_biwt, var_output_rsci_bdwt, var_output_rsci_bcwt, var_output_rsci_ivld_core_sct
);
  input core_wen;
  input var_output_rsci_oswt_unreg;
  input var_output_rsci_iswt0;
  input var_output_rsci_irdy;
  output var_output_rsci_biwt;
  output var_output_rsci_bdwt;
  input var_output_rsci_bcwt;
  output var_output_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire var_output_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign var_output_rsci_bdwt = var_output_rsci_oswt_unreg & core_wen;
  assign var_output_rsci_biwt = var_output_rsci_ogwt & var_output_rsci_irdy;
  assign var_output_rsci_ogwt = var_output_rsci_iswt0 & (~ var_output_rsci_bcwt);
  assign var_output_rsci_ivld_core_sct = var_output_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci_plm_kernel_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci_plm_kernel_wait_dp
    (
  clk, rst, plm_kernel_rsci_oswt_unreg, plm_kernel_rsci_bawt, plm_kernel_rsci_wen_comp,
      plm_kernel_rsci_idat_mxwt, plm_kernel_rsci_biwt, plm_kernel_rsci_bdwt, plm_kernel_rsci_bcwt,
      plm_kernel_rsci_idat
);
  input clk;
  input rst;
  input plm_kernel_rsci_oswt_unreg;
  output plm_kernel_rsci_bawt;
  output plm_kernel_rsci_wen_comp;
  output [1567:0] plm_kernel_rsci_idat_mxwt;
  input plm_kernel_rsci_biwt;
  input plm_kernel_rsci_bdwt;
  output plm_kernel_rsci_bcwt;
  reg plm_kernel_rsci_bcwt;
  input [1567:0] plm_kernel_rsci_idat;


  // Interconnect Declarations
  reg [1567:0] plm_kernel_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_kernel_rsci_bawt = plm_kernel_rsci_biwt | plm_kernel_rsci_bcwt;
  assign plm_kernel_rsci_wen_comp = (~ plm_kernel_rsci_oswt_unreg) | plm_kernel_rsci_bawt;
  assign plm_kernel_rsci_idat_mxwt = MUX_v_1568_2_2(plm_kernel_rsci_idat, plm_kernel_rsci_idat_bfwt,
      plm_kernel_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_kernel_rsci_bcwt <= ~((~(plm_kernel_rsci_bcwt | plm_kernel_rsci_biwt))
          | plm_kernel_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_bfwt <= {784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( plm_kernel_rsci_biwt ) begin
      plm_kernel_rsci_idat_bfwt <= plm_kernel_rsci_idat;
    end
  end

  function automatic [1567:0] MUX_v_1568_2_2;
    input [1567:0] input_0;
    input [1567:0] input_1;
    input [0:0] sel;
    reg [1567:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_1568_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci_plm_kernel_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci_plm_kernel_wait_ctrl
    (
  core_wen, plm_kernel_rsci_oswt_unreg, plm_kernel_rsci_iswt0, plm_kernel_rsci_biwt,
      plm_kernel_rsci_bdwt, plm_kernel_rsci_bcwt, plm_kernel_rsci_irdy_core_sct,
      plm_kernel_rsci_ivld
);
  input core_wen;
  input plm_kernel_rsci_oswt_unreg;
  input plm_kernel_rsci_iswt0;
  output plm_kernel_rsci_biwt;
  output plm_kernel_rsci_bdwt;
  input plm_kernel_rsci_bcwt;
  output plm_kernel_rsci_irdy_core_sct;
  input plm_kernel_rsci_ivld;


  // Interconnect Declarations
  wire plm_kernel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_kernel_rsci_bdwt = plm_kernel_rsci_oswt_unreg & core_wen;
  assign plm_kernel_rsci_biwt = plm_kernel_rsci_ogwt & plm_kernel_rsci_ivld;
  assign plm_kernel_rsci_ogwt = plm_kernel_rsci_iswt0 & (~ plm_kernel_rsci_bcwt);
  assign plm_kernel_rsci_irdy_core_sct = plm_kernel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci_buf_linear_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci_buf_linear_wait_dp
    (
  clk, rst, buf_linear_rsci_oswt_unreg, buf_linear_rsci_bawt, buf_linear_rsci_wen_comp,
      buf_linear_rsci_idat_mxwt, buf_linear_rsci_biwt, buf_linear_rsci_bdwt, buf_linear_rsci_bcwt,
      buf_linear_rsci_idat
);
  input clk;
  input rst;
  input buf_linear_rsci_oswt_unreg;
  output buf_linear_rsci_bawt;
  output buf_linear_rsci_wen_comp;
  output [4031:0] buf_linear_rsci_idat_mxwt;
  input buf_linear_rsci_biwt;
  input buf_linear_rsci_bdwt;
  output buf_linear_rsci_bcwt;
  reg buf_linear_rsci_bcwt;
  input [4031:0] buf_linear_rsci_idat;


  // Interconnect Declarations
  reg [4031:0] buf_linear_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign buf_linear_rsci_bawt = buf_linear_rsci_biwt | buf_linear_rsci_bcwt;
  assign buf_linear_rsci_wen_comp = (~ buf_linear_rsci_oswt_unreg) | buf_linear_rsci_bawt;
  assign buf_linear_rsci_idat_mxwt = MUX_v_4032_2_2(buf_linear_rsci_idat, buf_linear_rsci_idat_bfwt,
      buf_linear_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_bcwt <= 1'b0;
    end
    else begin
      buf_linear_rsci_bcwt <= ~((~(buf_linear_rsci_bcwt | buf_linear_rsci_biwt))
          | buf_linear_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_bfwt <= {504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( buf_linear_rsci_biwt ) begin
      buf_linear_rsci_idat_bfwt <= buf_linear_rsci_idat;
    end
  end

  function automatic [4031:0] MUX_v_4032_2_2;
    input [4031:0] input_0;
    input [4031:0] input_1;
    input [0:0] sel;
    reg [4031:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4032_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci_buf_linear_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci_buf_linear_wait_ctrl
    (
  core_wen, buf_linear_rsci_oswt_unreg, buf_linear_rsci_iswt0, buf_linear_rsci_biwt,
      buf_linear_rsci_bdwt, buf_linear_rsci_bcwt, buf_linear_rsci_irdy_core_sct,
      buf_linear_rsci_ivld
);
  input core_wen;
  input buf_linear_rsci_oswt_unreg;
  input buf_linear_rsci_iswt0;
  output buf_linear_rsci_biwt;
  output buf_linear_rsci_bdwt;
  input buf_linear_rsci_bcwt;
  output buf_linear_rsci_irdy_core_sct;
  input buf_linear_rsci_ivld;


  // Interconnect Declarations
  wire buf_linear_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign buf_linear_rsci_bdwt = buf_linear_rsci_oswt_unreg & core_wen;
  assign buf_linear_rsci_biwt = buf_linear_rsci_ogwt & buf_linear_rsci_ivld;
  assign buf_linear_rsci_ogwt = buf_linear_rsci_iswt0 & (~ buf_linear_rsci_bcwt);
  assign buf_linear_rsci_irdy_core_sct = buf_linear_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_dp
    (
  clk, rst, conf_info_rsci_oswt_unreg, conf_info_rsci_bawt, conf_info_rsci_wen_comp,
      conf_info_rsci_idat_mxwt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  wire [231:0] conf_info_rsci_idat_mxwt_pconst;
  reg [231:0] conf_info_rsci_idat_bfwt_231_0;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bawt = conf_info_rsci_biwt | conf_info_rsci_bcwt;
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt_unreg) | conf_info_rsci_bawt;
  assign conf_info_rsci_idat_mxwt_pconst = MUX_v_232_2_2((conf_info_rsci_idat[231:0]),
      conf_info_rsci_idat_bfwt_231_0, conf_info_rsci_bcwt);
  assign conf_info_rsci_idat_mxwt = {(conf_info_rsci_idat_mxwt_pconst[231:224]) ,
      (conf_info_rsci_idat_mxwt_pconst[199:192]) , (conf_info_rsci_idat_mxwt_pconst[167:160])
      , (conf_info_rsci_idat_mxwt_pconst[135:128]) , (conf_info_rsci_idat_mxwt_pconst[103:96])
      , (conf_info_rsci_idat_mxwt_pconst[71:64]) , (conf_info_rsci_idat_mxwt_pconst[39:32])
      , (conf_info_rsci_idat_mxwt_pconst[7:0])};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt_231_0 <= conf_info_rsci_idat[231:0];
    end
  end

  function automatic [231:0] MUX_v_232_2_2;
    input [231:0] input_0;
    input [231:0] input_1;
    input [0:0] sel;
    reg [231:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_232_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt_unreg, conf_info_rsci_iswt0, conf_info_rsci_biwt,
      conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt_unreg & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_iswt0 & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2dlb_cxx_catapult_store_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2dlb_cxx_catapult_store_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_staller (
  core_wen, conf_info_rsci_wen_comp, var_output_rsci_wen_comp, dma_write_ctrl_rsci_wen_comp,
      dma_write_chnl_rsci_wen_comp, done_rsci_wen_comp
);
  output core_wen;
  input conf_info_rsci_wen_comp;
  input var_output_rsci_wen_comp;
  input dma_write_ctrl_rsci_wen_comp;
  input dma_write_chnl_rsci_wen_comp;
  input done_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & var_output_rsci_wen_comp & dma_write_ctrl_rsci_wen_comp
      & dma_write_chnl_rsci_wen_comp & done_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt_unreg, done_rsci_bawt, done_rsci_wen_comp, done_rsci_biwt,
      done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bawt = done_rsci_biwt | done_rsci_bcwt;
  assign done_rsci_wen_comp = (~ done_rsci_oswt_unreg) | done_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt_unreg, done_rsci_iswt0, done_rsci_biwt, done_rsci_bdwt,
      done_rsci_bcwt, done_rsci_ivld_core_sct, done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt_unreg;
  input done_rsci_iswt0;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt_unreg & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_iswt0 & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
    (
  clk, rst, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_bawt, dma_write_chnl_rsci_wen_comp,
      dma_write_chnl_rsci_biwt, dma_write_chnl_rsci_bdwt, dma_write_chnl_rsci_bcwt
);
  input clk;
  input rst;
  input dma_write_chnl_rsci_oswt_unreg;
  output dma_write_chnl_rsci_bawt;
  output dma_write_chnl_rsci_wen_comp;
  input dma_write_chnl_rsci_biwt;
  input dma_write_chnl_rsci_bdwt;
  output dma_write_chnl_rsci_bcwt;
  reg dma_write_chnl_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_rsci_bawt = dma_write_chnl_rsci_biwt | dma_write_chnl_rsci_bcwt;
  assign dma_write_chnl_rsci_wen_comp = (~ dma_write_chnl_rsci_oswt_unreg) | dma_write_chnl_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_write_chnl_rsci_bcwt <= ~((~(dma_write_chnl_rsci_bcwt | dma_write_chnl_rsci_biwt))
          | dma_write_chnl_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
    (
  core_wen, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_iswt0, dma_write_chnl_rsci_irdy,
      dma_write_chnl_rsci_biwt, dma_write_chnl_rsci_bdwt, dma_write_chnl_rsci_bcwt,
      dma_write_chnl_rsci_ivld_core_sct
);
  input core_wen;
  input dma_write_chnl_rsci_oswt_unreg;
  input dma_write_chnl_rsci_iswt0;
  input dma_write_chnl_rsci_irdy;
  output dma_write_chnl_rsci_biwt;
  output dma_write_chnl_rsci_bdwt;
  input dma_write_chnl_rsci_bcwt;
  output dma_write_chnl_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire dma_write_chnl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_rsci_bdwt = dma_write_chnl_rsci_oswt_unreg & core_wen;
  assign dma_write_chnl_rsci_biwt = dma_write_chnl_rsci_ogwt & dma_write_chnl_rsci_irdy;
  assign dma_write_chnl_rsci_ogwt = dma_write_chnl_rsci_iswt0 & (~ dma_write_chnl_rsci_bcwt);
  assign dma_write_chnl_rsci_ivld_core_sct = dma_write_chnl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
    (
  clk, rst, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_bawt, dma_write_ctrl_rsci_wen_comp,
      dma_write_ctrl_rsci_biwt, dma_write_ctrl_rsci_bdwt, dma_write_ctrl_rsci_bcwt
);
  input clk;
  input rst;
  input dma_write_ctrl_rsci_oswt_unreg;
  output dma_write_ctrl_rsci_bawt;
  output dma_write_ctrl_rsci_wen_comp;
  input dma_write_ctrl_rsci_biwt;
  input dma_write_ctrl_rsci_bdwt;
  output dma_write_ctrl_rsci_bcwt;
  reg dma_write_ctrl_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_rsci_bawt = dma_write_ctrl_rsci_biwt | dma_write_ctrl_rsci_bcwt;
  assign dma_write_ctrl_rsci_wen_comp = (~ dma_write_ctrl_rsci_oswt_unreg) | dma_write_ctrl_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_rsci_bcwt <= ~((~(dma_write_ctrl_rsci_bcwt | dma_write_ctrl_rsci_biwt))
          | dma_write_ctrl_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
    (
  core_wen, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_iswt0, dma_write_ctrl_rsci_irdy,
      dma_write_ctrl_rsci_biwt, dma_write_ctrl_rsci_bdwt, dma_write_ctrl_rsci_bcwt,
      dma_write_ctrl_rsci_ivld_core_sct
);
  input core_wen;
  input dma_write_ctrl_rsci_oswt_unreg;
  input dma_write_ctrl_rsci_iswt0;
  input dma_write_ctrl_rsci_irdy;
  output dma_write_ctrl_rsci_biwt;
  output dma_write_ctrl_rsci_bdwt;
  input dma_write_ctrl_rsci_bcwt;
  output dma_write_ctrl_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire dma_write_ctrl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_rsci_bdwt = dma_write_ctrl_rsci_oswt_unreg & core_wen;
  assign dma_write_ctrl_rsci_biwt = dma_write_ctrl_rsci_ogwt & dma_write_ctrl_rsci_irdy;
  assign dma_write_ctrl_rsci_ogwt = dma_write_ctrl_rsci_iswt0 & (~ dma_write_ctrl_rsci_bcwt);
  assign dma_write_ctrl_rsci_ivld_core_sct = dma_write_ctrl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci_var_output_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci_var_output_wait_dp
    (
  clk, rst, var_output_rsci_oswt_unreg, var_output_rsci_bawt, var_output_rsci_wen_comp,
      var_output_rsci_idat_mxwt, var_output_rsci_biwt, var_output_rsci_bdwt, var_output_rsci_bcwt,
      var_output_rsci_idat
);
  input clk;
  input rst;
  input var_output_rsci_oswt_unreg;
  output var_output_rsci_bawt;
  output var_output_rsci_wen_comp;
  output [31:0] var_output_rsci_idat_mxwt;
  input var_output_rsci_biwt;
  input var_output_rsci_bdwt;
  output var_output_rsci_bcwt;
  reg var_output_rsci_bcwt;
  input [31:0] var_output_rsci_idat;


  // Interconnect Declarations
  reg [31:0] var_output_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign var_output_rsci_bawt = var_output_rsci_biwt | var_output_rsci_bcwt;
  assign var_output_rsci_wen_comp = (~ var_output_rsci_oswt_unreg) | var_output_rsci_bawt;
  assign var_output_rsci_idat_mxwt = MUX_v_32_2_2(var_output_rsci_idat, var_output_rsci_idat_bfwt,
      var_output_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      var_output_rsci_bcwt <= 1'b0;
    end
    else begin
      var_output_rsci_bcwt <= ~((~(var_output_rsci_bcwt | var_output_rsci_biwt))
          | var_output_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      var_output_rsci_idat_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( var_output_rsci_biwt ) begin
      var_output_rsci_idat_bfwt <= var_output_rsci_idat;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci_var_output_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci_var_output_wait_ctrl
    (
  core_wen, var_output_rsci_oswt_unreg, var_output_rsci_iswt0, var_output_rsci_biwt,
      var_output_rsci_bdwt, var_output_rsci_bcwt, var_output_rsci_irdy_core_sct,
      var_output_rsci_ivld
);
  input core_wen;
  input var_output_rsci_oswt_unreg;
  input var_output_rsci_iswt0;
  output var_output_rsci_biwt;
  output var_output_rsci_bdwt;
  input var_output_rsci_bcwt;
  output var_output_rsci_irdy_core_sct;
  input var_output_rsci_ivld;


  // Interconnect Declarations
  wire var_output_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign var_output_rsci_bdwt = var_output_rsci_oswt_unreg & core_wen;
  assign var_output_rsci_biwt = var_output_rsci_ogwt & var_output_rsci_ivld;
  assign var_output_rsci_ogwt = var_output_rsci_iswt0 & (~ var_output_rsci_bcwt);
  assign var_output_rsci_irdy_core_sct = var_output_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_dp
    (
  clk, rst, conf_info_rsci_oswt_unreg, conf_info_rsci_bawt, conf_info_rsci_wen_comp,
      conf_info_rsci_idat_mxwt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  wire [231:0] conf_info_rsci_idat_mxwt_pconst;
  reg [231:0] conf_info_rsci_idat_bfwt_231_0;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bawt = conf_info_rsci_biwt | conf_info_rsci_bcwt;
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt_unreg) | conf_info_rsci_bawt;
  assign conf_info_rsci_idat_mxwt_pconst = MUX_v_232_2_2((conf_info_rsci_idat[231:0]),
      conf_info_rsci_idat_bfwt_231_0, conf_info_rsci_bcwt);
  assign conf_info_rsci_idat_mxwt = {(conf_info_rsci_idat_mxwt_pconst[231:224]) ,
      (conf_info_rsci_idat_mxwt_pconst[199:192]) , (conf_info_rsci_idat_mxwt_pconst[167:160])
      , (conf_info_rsci_idat_mxwt_pconst[135:128]) , (conf_info_rsci_idat_mxwt_pconst[103:96])
      , (conf_info_rsci_idat_mxwt_pconst[71:64]) , (conf_info_rsci_idat_mxwt_pconst[39:32])
      , (conf_info_rsci_idat_mxwt_pconst[7:0])};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt_231_0 <= conf_info_rsci_idat[231:0];
    end
  end

  function automatic [231:0] MUX_v_232_2_2;
    input [231:0] input_0;
    input [231:0] input_1;
    input [0:0] sel;
    reg [231:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_232_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt_unreg, conf_info_rsci_iswt0, conf_info_rsci_biwt,
      conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt_unreg & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_iswt0 & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi
    (
  clk, rst, store_done_cns_rdy, store_done_cns_vld, core_wen, store_done_cnsi_oswt_unreg,
      store_done_cnsi_bawt, store_done_cnsi_iswt0, store_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output store_done_cns_rdy;
  input store_done_cns_vld;
  input core_wen;
  input store_done_cnsi_oswt_unreg;
  output store_done_cnsi_bawt;
  input store_done_cnsi_iswt0;
  output store_done_cnsi_wen_comp;


  // Interconnect Declarations
  wire store_done_cnsi_ivld;
  wire store_done_cnsi_biwt;
  wire store_done_cnsi_bdwt;
  wire store_done_cnsi_bcwt;
  wire store_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd48)) store_done_cnsi
      (
      .vld(store_done_cns_vld),
      .rdy(store_done_cns_rdy),
      .ivld(store_done_cnsi_ivld),
      .irdy(store_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl
      conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl_inst (
      .core_wen(core_wen),
      .store_done_cnsi_oswt_unreg(store_done_cnsi_oswt_unreg),
      .store_done_cnsi_iswt0(store_done_cnsi_iswt0),
      .store_done_cnsi_ivld(store_done_cnsi_ivld),
      .store_done_cnsi_biwt(store_done_cnsi_biwt),
      .store_done_cnsi_bdwt(store_done_cnsi_bdwt),
      .store_done_cnsi_bcwt(store_done_cnsi_bcwt),
      .store_done_cnsi_irdy_core_sct(store_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp
      conv2dlb_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .store_done_cnsi_oswt_unreg(store_done_cnsi_oswt_unreg),
      .store_done_cnsi_bawt(store_done_cnsi_bawt),
      .store_done_cnsi_wen_comp(store_done_cnsi_wen_comp),
      .store_done_cnsi_biwt(store_done_cnsi_biwt),
      .store_done_cnsi_bdwt(store_done_cnsi_bdwt),
      .store_done_cnsi_bcwt(store_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi
    (
  clk, rst, compute_done_cns_rdy, compute_done_cns_vld, core_wen, compute_done_cnsi_oswt_unreg,
      compute_done_cnsi_bawt, compute_done_cnsi_iswt0, compute_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output compute_done_cns_rdy;
  input compute_done_cns_vld;
  input core_wen;
  input compute_done_cnsi_oswt_unreg;
  output compute_done_cnsi_bawt;
  input compute_done_cnsi_iswt0;
  output compute_done_cnsi_wen_comp;


  // Interconnect Declarations
  wire compute_done_cnsi_ivld;
  wire compute_done_cnsi_biwt;
  wire compute_done_cnsi_bdwt;
  wire compute_done_cnsi_bcwt;
  wire compute_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd47)) compute_done_cnsi
      (
      .vld(compute_done_cns_vld),
      .rdy(compute_done_cns_rdy),
      .ivld(compute_done_cnsi_ivld),
      .irdy(compute_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl
      conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .compute_done_cnsi_oswt_unreg(compute_done_cnsi_oswt_unreg),
      .compute_done_cnsi_iswt0(compute_done_cnsi_iswt0),
      .compute_done_cnsi_ivld(compute_done_cnsi_ivld),
      .compute_done_cnsi_biwt(compute_done_cnsi_biwt),
      .compute_done_cnsi_bdwt(compute_done_cnsi_bdwt),
      .compute_done_cnsi_bcwt(compute_done_cnsi_bcwt),
      .compute_done_cnsi_irdy_core_sct(compute_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp
      conv2dlb_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_done_cnsi_oswt_unreg(compute_done_cnsi_oswt_unreg),
      .compute_done_cnsi_bawt(compute_done_cnsi_bawt),
      .compute_done_cnsi_wen_comp(compute_done_cnsi_wen_comp),
      .compute_done_cnsi_biwt(compute_done_cnsi_biwt),
      .compute_done_cnsi_bdwt(compute_done_cnsi_bdwt),
      .compute_done_cnsi_bcwt(compute_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi
    (
  clk, rst, load_done_cns_rdy, load_done_cns_vld, core_wen, load_done_cnsi_oswt_unreg,
      load_done_cnsi_bawt, load_done_cnsi_iswt0, load_done_cnsi_wen_comp, load_done_cnsi_irdy_core_psct
);
  input clk;
  input rst;
  output load_done_cns_rdy;
  input load_done_cns_vld;
  input core_wen;
  input load_done_cnsi_oswt_unreg;
  output load_done_cnsi_bawt;
  input load_done_cnsi_iswt0;
  output load_done_cnsi_wen_comp;
  input load_done_cnsi_irdy_core_psct;


  // Interconnect Declarations
  wire load_done_cnsi_ivld;
  wire load_done_cnsi_biwt;
  wire load_done_cnsi_bdwt;
  wire load_done_cnsi_bcwt;
  wire load_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd46)) load_done_cnsi
      (
      .vld(load_done_cns_vld),
      .rdy(load_done_cns_rdy),
      .ivld(load_done_cnsi_ivld),
      .irdy(load_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl
      conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl_inst (
      .core_wen(core_wen),
      .load_done_cnsi_oswt_unreg(load_done_cnsi_oswt_unreg),
      .load_done_cnsi_iswt0(load_done_cnsi_iswt0),
      .load_done_cnsi_irdy_core_psct(load_done_cnsi_irdy_core_psct),
      .load_done_cnsi_ivld(load_done_cnsi_ivld),
      .load_done_cnsi_biwt(load_done_cnsi_biwt),
      .load_done_cnsi_bdwt(load_done_cnsi_bdwt),
      .load_done_cnsi_bcwt(load_done_cnsi_bcwt),
      .load_done_cnsi_irdy_core_sct(load_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp
      conv2dlb_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .load_done_cnsi_oswt_unreg(load_done_cnsi_oswt_unreg),
      .load_done_cnsi_bawt(load_done_cnsi_bawt),
      .load_done_cnsi_wen_comp(load_done_cnsi_wen_comp),
      .load_done_cnsi_biwt(load_done_cnsi_biwt),
      .load_done_cnsi_bdwt(load_done_cnsi_bdwt),
      .load_done_cnsi_bcwt(load_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi
    (
  clk, rst, config_done_cns_rdy, config_done_cns_vld, core_wen, config_done_cnsi_oswt_unreg,
      config_done_cnsi_bawt, config_done_cnsi_iswt0, config_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output config_done_cns_rdy;
  input config_done_cns_vld;
  input core_wen;
  input config_done_cnsi_oswt_unreg;
  output config_done_cnsi_bawt;
  input config_done_cnsi_iswt0;
  output config_done_cnsi_wen_comp;


  // Interconnect Declarations
  wire config_done_cnsi_ivld;
  wire config_done_cnsi_biwt;
  wire config_done_cnsi_bdwt;
  wire config_done_cnsi_bcwt;
  wire config_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd45)) config_done_cnsi
      (
      .vld(config_done_cns_vld),
      .rdy(config_done_cns_rdy),
      .ivld(config_done_cnsi_ivld),
      .irdy(config_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl
      conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .config_done_cnsi_oswt_unreg(config_done_cnsi_oswt_unreg),
      .config_done_cnsi_iswt0(config_done_cnsi_iswt0),
      .config_done_cnsi_ivld(config_done_cnsi_ivld),
      .config_done_cnsi_biwt(config_done_cnsi_biwt),
      .config_done_cnsi_bdwt(config_done_cnsi_bdwt),
      .config_done_cnsi_bcwt(config_done_cnsi_bcwt),
      .config_done_cnsi_irdy_core_sct(config_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp
      conv2dlb_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .config_done_cnsi_oswt_unreg(config_done_cnsi_oswt_unreg),
      .config_done_cnsi_bawt(config_done_cnsi_bawt),
      .config_done_cnsi_wen_comp(config_done_cnsi_wen_comp),
      .config_done_cnsi_biwt(config_done_cnsi_biwt),
      .config_done_cnsi_bdwt(config_done_cnsi_bdwt),
      .config_done_cnsi_bcwt(config_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci
    (
  clk, rst, acc_done_rsc_vld, core_wen, acc_done_rsci_oswt_unreg, acc_done_rsci_bawt,
      acc_done_rsci_iswt0, core_wten
);
  input clk;
  input rst;
  output acc_done_rsc_vld;
  input core_wen;
  input acc_done_rsci_oswt_unreg;
  output acc_done_rsci_bawt;
  input acc_done_rsci_iswt0;
  input core_wten;


  // Interconnect Declarations
  wire acc_done_rsci_biwt;
  wire acc_done_rsci_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_out_vld_v1 #(.rscid(32'sd44)) acc_done_rsci
      (
      .vld(acc_done_rsc_vld),
      .ivld(acc_done_rsci_biwt)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl
      conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl_inst (
      .core_wen(core_wen),
      .acc_done_rsci_oswt_unreg(acc_done_rsci_oswt_unreg),
      .acc_done_rsci_iswt0(acc_done_rsci_iswt0),
      .core_wten(core_wten),
      .acc_done_rsci_biwt(acc_done_rsci_biwt),
      .acc_done_rsci_bdwt(acc_done_rsci_bdwt)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp
      conv2dlb_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .acc_done_rsci_bawt(acc_done_rsci_bawt),
      .acc_done_rsci_biwt(acc_done_rsci_biwt),
      .acc_done_rsci_bdwt(acc_done_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt_unreg, done_rsci_bawt,
      done_rsci_iswt0, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  input done_rsci_iswt0;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd5)) done_rsci
      (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci_done_wait_ctrl config_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_iswt0(done_rsci_iswt0),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci_done_wait_dp config_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci (
  clk, rst, plm_conf_store_rsc_dat, plm_conf_store_rsc_vld, plm_conf_store_rsc_rdy,
      core_wen, plm_conf_store_rsci_oswt_unreg, plm_conf_store_rsci_bawt, plm_conf_store_rsci_iswt0,
      plm_conf_store_rsci_wen_comp, plm_conf_store_rsci_idat
);
  input clk;
  input rst;
  output [255:0] plm_conf_store_rsc_dat;
  output plm_conf_store_rsc_vld;
  input plm_conf_store_rsc_rdy;
  input core_wen;
  input plm_conf_store_rsci_oswt_unreg;
  output plm_conf_store_rsci_bawt;
  input plm_conf_store_rsci_iswt0;
  output plm_conf_store_rsci_wen_comp;
  input [255:0] plm_conf_store_rsci_idat;


  // Interconnect Declarations
  wire plm_conf_store_rsci_irdy;
  wire plm_conf_store_rsci_biwt;
  wire plm_conf_store_rsci_bdwt;
  wire plm_conf_store_rsci_bcwt;
  wire plm_conf_store_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd256)) plm_conf_store_rsci (
      .irdy(plm_conf_store_rsci_irdy),
      .ivld(plm_conf_store_rsci_ivld_core_sct),
      .idat(plm_conf_store_rsci_idat),
      .rdy(plm_conf_store_rsc_rdy),
      .vld(plm_conf_store_rsc_vld),
      .dat(plm_conf_store_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl
      config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_conf_store_rsci_oswt_unreg(plm_conf_store_rsci_oswt_unreg),
      .plm_conf_store_rsci_iswt0(plm_conf_store_rsci_iswt0),
      .plm_conf_store_rsci_irdy(plm_conf_store_rsci_irdy),
      .plm_conf_store_rsci_biwt(plm_conf_store_rsci_biwt),
      .plm_conf_store_rsci_bdwt(plm_conf_store_rsci_bdwt),
      .plm_conf_store_rsci_bcwt(plm_conf_store_rsci_bcwt),
      .plm_conf_store_rsci_ivld_core_sct(plm_conf_store_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_dp
      config_core_plm_conf_store_rsci_plm_conf_store_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_conf_store_rsci_oswt_unreg(plm_conf_store_rsci_oswt_unreg),
      .plm_conf_store_rsci_bawt(plm_conf_store_rsci_bawt),
      .plm_conf_store_rsci_wen_comp(plm_conf_store_rsci_wen_comp),
      .plm_conf_store_rsci_biwt(plm_conf_store_rsci_biwt),
      .plm_conf_store_rsci_bdwt(plm_conf_store_rsci_bdwt),
      .plm_conf_store_rsci_bcwt(plm_conf_store_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci (
  clk, rst, plm_conf_compute_rsc_dat, plm_conf_compute_rsc_vld, plm_conf_compute_rsc_rdy,
      core_wen, plm_conf_compute_rsci_oswt_unreg, plm_conf_compute_rsci_bawt, plm_conf_compute_rsci_iswt0,
      plm_conf_compute_rsci_wen_comp, plm_conf_compute_rsci_idat
);
  input clk;
  input rst;
  output [255:0] plm_conf_compute_rsc_dat;
  output plm_conf_compute_rsc_vld;
  input plm_conf_compute_rsc_rdy;
  input core_wen;
  input plm_conf_compute_rsci_oswt_unreg;
  output plm_conf_compute_rsci_bawt;
  input plm_conf_compute_rsci_iswt0;
  output plm_conf_compute_rsci_wen_comp;
  input [255:0] plm_conf_compute_rsci_idat;


  // Interconnect Declarations
  wire plm_conf_compute_rsci_irdy;
  wire plm_conf_compute_rsci_biwt;
  wire plm_conf_compute_rsci_bdwt;
  wire plm_conf_compute_rsci_bcwt;
  wire plm_conf_compute_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd256)) plm_conf_compute_rsci (
      .irdy(plm_conf_compute_rsci_irdy),
      .ivld(plm_conf_compute_rsci_ivld_core_sct),
      .idat(plm_conf_compute_rsci_idat),
      .rdy(plm_conf_compute_rsc_rdy),
      .vld(plm_conf_compute_rsc_vld),
      .dat(plm_conf_compute_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl
      config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_conf_compute_rsci_oswt_unreg(plm_conf_compute_rsci_oswt_unreg),
      .plm_conf_compute_rsci_iswt0(plm_conf_compute_rsci_iswt0),
      .plm_conf_compute_rsci_irdy(plm_conf_compute_rsci_irdy),
      .plm_conf_compute_rsci_biwt(plm_conf_compute_rsci_biwt),
      .plm_conf_compute_rsci_bdwt(plm_conf_compute_rsci_bdwt),
      .plm_conf_compute_rsci_bcwt(plm_conf_compute_rsci_bcwt),
      .plm_conf_compute_rsci_ivld_core_sct(plm_conf_compute_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp
      config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_conf_compute_rsci_oswt_unreg(plm_conf_compute_rsci_oswt_unreg),
      .plm_conf_compute_rsci_bawt(plm_conf_compute_rsci_bawt),
      .plm_conf_compute_rsci_wen_comp(plm_conf_compute_rsci_wen_comp),
      .plm_conf_compute_rsci_biwt(plm_conf_compute_rsci_biwt),
      .plm_conf_compute_rsci_bdwt(plm_conf_compute_rsci_bdwt),
      .plm_conf_compute_rsci_bcwt(plm_conf_compute_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci (
  clk, rst, plm_conf_load_rsc_dat, plm_conf_load_rsc_vld, plm_conf_load_rsc_rdy,
      core_wen, plm_conf_load_rsci_oswt_unreg, plm_conf_load_rsci_bawt, plm_conf_load_rsci_iswt0,
      plm_conf_load_rsci_wen_comp, plm_conf_load_rsci_idat
);
  input clk;
  input rst;
  output [255:0] plm_conf_load_rsc_dat;
  output plm_conf_load_rsc_vld;
  input plm_conf_load_rsc_rdy;
  input core_wen;
  input plm_conf_load_rsci_oswt_unreg;
  output plm_conf_load_rsci_bawt;
  input plm_conf_load_rsci_iswt0;
  output plm_conf_load_rsci_wen_comp;
  input [255:0] plm_conf_load_rsci_idat;


  // Interconnect Declarations
  wire plm_conf_load_rsci_irdy;
  wire plm_conf_load_rsci_biwt;
  wire plm_conf_load_rsci_bdwt;
  wire plm_conf_load_rsci_bcwt;
  wire plm_conf_load_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd256)) plm_conf_load_rsci (
      .irdy(plm_conf_load_rsci_irdy),
      .ivld(plm_conf_load_rsci_ivld_core_sct),
      .idat(plm_conf_load_rsci_idat),
      .rdy(plm_conf_load_rsc_rdy),
      .vld(plm_conf_load_rsc_vld),
      .dat(plm_conf_load_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl
      config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_conf_load_rsci_oswt_unreg(plm_conf_load_rsci_oswt_unreg),
      .plm_conf_load_rsci_iswt0(plm_conf_load_rsci_iswt0),
      .plm_conf_load_rsci_irdy(plm_conf_load_rsci_irdy),
      .plm_conf_load_rsci_biwt(plm_conf_load_rsci_biwt),
      .plm_conf_load_rsci_bdwt(plm_conf_load_rsci_bdwt),
      .plm_conf_load_rsci_bcwt(plm_conf_load_rsci_bcwt),
      .plm_conf_load_rsci_ivld_core_sct(plm_conf_load_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_dp
      config_core_plm_conf_load_rsci_plm_conf_load_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_conf_load_rsci_oswt_unreg(plm_conf_load_rsci_oswt_unreg),
      .plm_conf_load_rsci_bawt(plm_conf_load_rsci_bawt),
      .plm_conf_load_rsci_wen_comp(plm_conf_load_rsci_wen_comp),
      .plm_conf_load_rsci_biwt(plm_conf_load_rsci_biwt),
      .plm_conf_load_rsci_bdwt(plm_conf_load_rsci_bdwt),
      .plm_conf_load_rsci_bcwt(plm_conf_load_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt_unreg,
      conf_info_rsci_bawt, conf_info_rsci_iswt0, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_wen_comp;
  output [255:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_ctrl config_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_iswt0(conf_info_rsci_iswt0),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_dp config_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1
    (
  clk, rst, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  input [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1;
  output [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff;
  input LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_ctrl
      load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_core_sct_pff(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_core_sct_iff),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_dp
      load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_biwt_1),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bdwt_2)
    );
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff = LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_core_sct_iff;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d =
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd11)) done_rsci
      (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci_done_wait_ctrl load_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt(done_rsci_oswt),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci_done_wait_dp load_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt(done_rsci_oswt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci (
  clk, rst, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy,
      core_wen, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_bawt, dma_read_chnl_rsci_iswt0,
      dma_read_chnl_rsci_wen_comp, dma_read_chnl_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  input core_wen;
  input dma_read_chnl_rsci_oswt_unreg;
  output dma_read_chnl_rsci_bawt;
  input dma_read_chnl_rsci_iswt0;
  output dma_read_chnl_rsci_wen_comp;
  output [31:0] dma_read_chnl_rsci_idat_mxwt;


  // Interconnect Declarations
  wire dma_read_chnl_rsci_biwt;
  wire dma_read_chnl_rsci_bdwt;
  wire dma_read_chnl_rsci_bcwt;
  wire dma_read_chnl_rsci_irdy_core_sct;
  wire dma_read_chnl_rsci_ivld;
  wire [63:0] dma_read_chnl_rsci_idat;
  wire [31:0] dma_read_chnl_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd10),
  .width(32'sd64)) dma_read_chnl_rsci (
      .rdy(dma_read_chnl_rsc_rdy),
      .vld(dma_read_chnl_rsc_vld),
      .dat(dma_read_chnl_rsc_dat),
      .irdy(dma_read_chnl_rsci_irdy_core_sct),
      .ivld(dma_read_chnl_rsci_ivld),
      .idat(dma_read_chnl_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
      load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl_inst (
      .core_wen(core_wen),
      .dma_read_chnl_rsci_oswt_unreg(dma_read_chnl_rsci_oswt_unreg),
      .dma_read_chnl_rsci_iswt0(dma_read_chnl_rsci_iswt0),
      .dma_read_chnl_rsci_biwt(dma_read_chnl_rsci_biwt),
      .dma_read_chnl_rsci_bdwt(dma_read_chnl_rsci_bdwt),
      .dma_read_chnl_rsci_bcwt(dma_read_chnl_rsci_bcwt),
      .dma_read_chnl_rsci_irdy_core_sct(dma_read_chnl_rsci_irdy_core_sct),
      .dma_read_chnl_rsci_ivld(dma_read_chnl_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
      load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_rsci_oswt_unreg(dma_read_chnl_rsci_oswt_unreg),
      .dma_read_chnl_rsci_bawt(dma_read_chnl_rsci_bawt),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .dma_read_chnl_rsci_idat_mxwt(dma_read_chnl_rsci_idat_mxwt_pconst),
      .dma_read_chnl_rsci_biwt(dma_read_chnl_rsci_biwt),
      .dma_read_chnl_rsci_bdwt(dma_read_chnl_rsci_bdwt),
      .dma_read_chnl_rsci_bcwt(dma_read_chnl_rsci_bcwt),
      .dma_read_chnl_rsci_idat(dma_read_chnl_rsci_idat)
    );
  assign dma_read_chnl_rsci_idat_mxwt = dma_read_chnl_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci (
  clk, rst, dma_read_ctrl_rsc_dat, dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy,
      core_wen, core_wten, dma_read_ctrl_rsci_oswt_unreg, dma_read_ctrl_rsci_bawt,
      dma_read_ctrl_rsci_iswt0, dma_read_ctrl_rsci_irdy_mxwt, dma_read_ctrl_rsci_idat
);
  input clk;
  input rst;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  input core_wen;
  input core_wten;
  input dma_read_ctrl_rsci_oswt_unreg;
  output dma_read_ctrl_rsci_bawt;
  input dma_read_ctrl_rsci_iswt0;
  output dma_read_ctrl_rsci_irdy_mxwt;
  input [66:0] dma_read_ctrl_rsci_idat;


  // Interconnect Declarations
  wire dma_read_ctrl_rsci_irdy;
  wire dma_read_ctrl_rsci_biwt;
  wire dma_read_ctrl_rsci_bdwt;


  // Interconnect Declarations for Component Instantiations 
  wire [66:0] nl_dma_read_ctrl_rsci_idat;
  assign nl_dma_read_ctrl_rsci_idat = {19'b0110000000000000000 , (dma_read_ctrl_rsci_idat[47:32])
      , 16'b0000000000000000 , (dma_read_ctrl_rsci_idat[15:0])};
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd9),
  .width(32'sd67)) dma_read_ctrl_rsci (
      .irdy(dma_read_ctrl_rsci_irdy),
      .ivld(dma_read_ctrl_rsci_biwt),
      .idat(nl_dma_read_ctrl_rsci_idat[66:0]),
      .rdy(dma_read_ctrl_rsc_rdy),
      .vld(dma_read_ctrl_rsc_vld),
      .dat(dma_read_ctrl_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
      load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dma_read_ctrl_rsci_oswt_unreg(dma_read_ctrl_rsci_oswt_unreg),
      .dma_read_ctrl_rsci_iswt0(dma_read_ctrl_rsci_iswt0),
      .dma_read_ctrl_rsci_biwt(dma_read_ctrl_rsci_biwt),
      .dma_read_ctrl_rsci_bdwt(dma_read_ctrl_rsci_bdwt)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
      load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_rsci_bawt(dma_read_ctrl_rsci_bawt),
      .dma_read_ctrl_rsci_irdy_mxwt(dma_read_ctrl_rsci_irdy_mxwt),
      .dma_read_ctrl_rsci_irdy(dma_read_ctrl_rsci_irdy),
      .dma_read_ctrl_rsci_biwt(dma_read_ctrl_rsci_biwt),
      .dma_read_ctrl_rsci_bdwt(dma_read_ctrl_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci (
  clk, rst, plm_kernel_rsc_dat, plm_kernel_rsc_vld, plm_kernel_rsc_rdy, core_wen,
      plm_kernel_rsci_oswt_unreg, plm_kernel_rsci_bawt, plm_kernel_rsci_iswt0, plm_kernel_rsci_wen_comp,
      plm_kernel_rsci_idat
);
  input clk;
  input rst;
  output [1567:0] plm_kernel_rsc_dat;
  output plm_kernel_rsc_vld;
  input plm_kernel_rsc_rdy;
  input core_wen;
  input plm_kernel_rsci_oswt_unreg;
  output plm_kernel_rsci_bawt;
  input plm_kernel_rsci_iswt0;
  output plm_kernel_rsci_wen_comp;
  input [1567:0] plm_kernel_rsci_idat;


  // Interconnect Declarations
  wire plm_kernel_rsci_irdy;
  wire plm_kernel_rsci_biwt;
  wire plm_kernel_rsci_bdwt;
  wire plm_kernel_rsci_bcwt;
  wire plm_kernel_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd8),
  .width(32'sd1568)) plm_kernel_rsci (
      .irdy(plm_kernel_rsci_irdy),
      .ivld(plm_kernel_rsci_ivld_core_sct),
      .idat(plm_kernel_rsci_idat),
      .rdy(plm_kernel_rsc_rdy),
      .vld(plm_kernel_rsc_vld),
      .dat(plm_kernel_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci_plm_kernel_wait_ctrl load_core_plm_kernel_rsci_plm_kernel_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .plm_kernel_rsci_oswt_unreg(plm_kernel_rsci_oswt_unreg),
      .plm_kernel_rsci_iswt0(plm_kernel_rsci_iswt0),
      .plm_kernel_rsci_irdy(plm_kernel_rsci_irdy),
      .plm_kernel_rsci_biwt(plm_kernel_rsci_biwt),
      .plm_kernel_rsci_bdwt(plm_kernel_rsci_bdwt),
      .plm_kernel_rsci_bcwt(plm_kernel_rsci_bcwt),
      .plm_kernel_rsci_ivld_core_sct(plm_kernel_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci_plm_kernel_wait_dp load_core_plm_kernel_rsci_plm_kernel_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_kernel_rsci_oswt_unreg(plm_kernel_rsci_oswt_unreg),
      .plm_kernel_rsci_bawt(plm_kernel_rsci_bawt),
      .plm_kernel_rsci_wen_comp(plm_kernel_rsci_wen_comp),
      .plm_kernel_rsci_biwt(plm_kernel_rsci_biwt),
      .plm_kernel_rsci_bdwt(plm_kernel_rsci_bdwt),
      .plm_kernel_rsci_bcwt(plm_kernel_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci (
  clk, rst, buf_linear_rsc_dat, buf_linear_rsc_vld, buf_linear_rsc_rdy, core_wen,
      buf_linear_rsci_oswt_unreg, buf_linear_rsci_bawt, buf_linear_rsci_iswt0, buf_linear_rsci_wen_comp,
      buf_linear_rsci_idat
);
  input clk;
  input rst;
  output [4031:0] buf_linear_rsc_dat;
  output buf_linear_rsc_vld;
  input buf_linear_rsc_rdy;
  input core_wen;
  input buf_linear_rsci_oswt_unreg;
  output buf_linear_rsci_bawt;
  input buf_linear_rsci_iswt0;
  output buf_linear_rsci_wen_comp;
  input [4031:0] buf_linear_rsci_idat;


  // Interconnect Declarations
  wire buf_linear_rsci_irdy;
  wire buf_linear_rsci_biwt;
  wire buf_linear_rsci_bdwt;
  wire buf_linear_rsci_bcwt;
  wire buf_linear_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd7),
  .width(32'sd4032)) buf_linear_rsci (
      .irdy(buf_linear_rsci_irdy),
      .ivld(buf_linear_rsci_ivld_core_sct),
      .idat(buf_linear_rsci_idat),
      .rdy(buf_linear_rsc_rdy),
      .vld(buf_linear_rsc_vld),
      .dat(buf_linear_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci_buf_linear_wait_ctrl load_core_buf_linear_rsci_buf_linear_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .buf_linear_rsci_oswt_unreg(buf_linear_rsci_oswt_unreg),
      .buf_linear_rsci_iswt0(buf_linear_rsci_iswt0),
      .buf_linear_rsci_irdy(buf_linear_rsci_irdy),
      .buf_linear_rsci_biwt(buf_linear_rsci_biwt),
      .buf_linear_rsci_bdwt(buf_linear_rsci_bdwt),
      .buf_linear_rsci_bcwt(buf_linear_rsci_bcwt),
      .buf_linear_rsci_ivld_core_sct(buf_linear_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci_buf_linear_wait_dp load_core_buf_linear_rsci_buf_linear_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .buf_linear_rsci_oswt_unreg(buf_linear_rsci_oswt_unreg),
      .buf_linear_rsci_bawt(buf_linear_rsci_bawt),
      .buf_linear_rsci_wen_comp(buf_linear_rsci_wen_comp),
      .buf_linear_rsci_biwt(buf_linear_rsci_biwt),
      .buf_linear_rsci_bdwt(buf_linear_rsci_bdwt),
      .buf_linear_rsci_bcwt(buf_linear_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt,
      conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt;
  output conf_info_rsci_wen_comp;
  output [231:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;
  wire [231:0] conf_info_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd6),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_ctrl load_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt(conf_info_rsci_oswt),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_dp load_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt(conf_info_rsci_oswt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt_pconst),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
  assign conf_info_rsci_idat_mxwt = conf_info_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt_unreg, done_rsci_bawt,
      done_rsci_iswt0, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  input done_rsci_iswt0;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd19)) done_rsci
      (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci_done_wait_ctrl compute_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_iswt0(done_rsci_iswt0),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci_done_wait_dp compute_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci (
  clk, rst, var_output_rsc_dat, var_output_rsc_vld, var_output_rsc_rdy, core_wen,
      var_output_rsci_oswt_unreg, var_output_rsci_bawt, var_output_rsci_iswt0, var_output_rsci_wen_comp,
      var_output_rsci_idat
);
  input clk;
  input rst;
  output [31:0] var_output_rsc_dat;
  output var_output_rsc_vld;
  input var_output_rsc_rdy;
  input core_wen;
  input var_output_rsci_oswt_unreg;
  output var_output_rsci_bawt;
  input var_output_rsci_iswt0;
  output var_output_rsci_wen_comp;
  input [31:0] var_output_rsci_idat;


  // Interconnect Declarations
  wire var_output_rsci_irdy;
  wire var_output_rsci_biwt;
  wire var_output_rsci_bdwt;
  wire var_output_rsci_bcwt;
  wire var_output_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd18),
  .width(32'sd32)) var_output_rsci (
      .irdy(var_output_rsci_irdy),
      .ivld(var_output_rsci_ivld_core_sct),
      .idat(var_output_rsci_idat),
      .rdy(var_output_rsc_rdy),
      .vld(var_output_rsc_vld),
      .dat(var_output_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci_var_output_wait_ctrl
      compute_core_var_output_rsci_var_output_wait_ctrl_inst (
      .core_wen(core_wen),
      .var_output_rsci_oswt_unreg(var_output_rsci_oswt_unreg),
      .var_output_rsci_iswt0(var_output_rsci_iswt0),
      .var_output_rsci_irdy(var_output_rsci_irdy),
      .var_output_rsci_biwt(var_output_rsci_biwt),
      .var_output_rsci_bdwt(var_output_rsci_bdwt),
      .var_output_rsci_bcwt(var_output_rsci_bcwt),
      .var_output_rsci_ivld_core_sct(var_output_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci_var_output_wait_dp compute_core_var_output_rsci_var_output_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .var_output_rsci_oswt_unreg(var_output_rsci_oswt_unreg),
      .var_output_rsci_bawt(var_output_rsci_bawt),
      .var_output_rsci_wen_comp(var_output_rsci_wen_comp),
      .var_output_rsci_biwt(var_output_rsci_biwt),
      .var_output_rsci_bdwt(var_output_rsci_bdwt),
      .var_output_rsci_bcwt(var_output_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci (
  clk, rst, plm_kernel_rsc_dat, plm_kernel_rsc_vld, plm_kernel_rsc_rdy, core_wen,
      plm_kernel_rsci_oswt_unreg, plm_kernel_rsci_bawt, plm_kernel_rsci_iswt0, plm_kernel_rsci_wen_comp,
      plm_kernel_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [1567:0] plm_kernel_rsc_dat;
  input plm_kernel_rsc_vld;
  output plm_kernel_rsc_rdy;
  input core_wen;
  input plm_kernel_rsci_oswt_unreg;
  output plm_kernel_rsci_bawt;
  input plm_kernel_rsci_iswt0;
  output plm_kernel_rsci_wen_comp;
  output [1567:0] plm_kernel_rsci_idat_mxwt;


  // Interconnect Declarations
  wire plm_kernel_rsci_biwt;
  wire plm_kernel_rsci_bdwt;
  wire plm_kernel_rsci_bcwt;
  wire plm_kernel_rsci_irdy_core_sct;
  wire plm_kernel_rsci_ivld;
  wire [1567:0] plm_kernel_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd17),
  .width(32'sd1568)) plm_kernel_rsci (
      .rdy(plm_kernel_rsc_rdy),
      .vld(plm_kernel_rsc_vld),
      .dat(plm_kernel_rsc_dat),
      .irdy(plm_kernel_rsci_irdy_core_sct),
      .ivld(plm_kernel_rsci_ivld),
      .idat(plm_kernel_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci_plm_kernel_wait_ctrl
      compute_core_plm_kernel_rsci_plm_kernel_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_kernel_rsci_oswt_unreg(plm_kernel_rsci_oswt_unreg),
      .plm_kernel_rsci_iswt0(plm_kernel_rsci_iswt0),
      .plm_kernel_rsci_biwt(plm_kernel_rsci_biwt),
      .plm_kernel_rsci_bdwt(plm_kernel_rsci_bdwt),
      .plm_kernel_rsci_bcwt(plm_kernel_rsci_bcwt),
      .plm_kernel_rsci_irdy_core_sct(plm_kernel_rsci_irdy_core_sct),
      .plm_kernel_rsci_ivld(plm_kernel_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci_plm_kernel_wait_dp compute_core_plm_kernel_rsci_plm_kernel_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_kernel_rsci_oswt_unreg(plm_kernel_rsci_oswt_unreg),
      .plm_kernel_rsci_bawt(plm_kernel_rsci_bawt),
      .plm_kernel_rsci_wen_comp(plm_kernel_rsci_wen_comp),
      .plm_kernel_rsci_idat_mxwt(plm_kernel_rsci_idat_mxwt),
      .plm_kernel_rsci_biwt(plm_kernel_rsci_biwt),
      .plm_kernel_rsci_bdwt(plm_kernel_rsci_bdwt),
      .plm_kernel_rsci_bcwt(plm_kernel_rsci_bcwt),
      .plm_kernel_rsci_idat(plm_kernel_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci (
  clk, rst, buf_linear_rsc_dat, buf_linear_rsc_vld, buf_linear_rsc_rdy, core_wen,
      buf_linear_rsci_oswt_unreg, buf_linear_rsci_bawt, buf_linear_rsci_iswt0, buf_linear_rsci_wen_comp,
      buf_linear_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [4031:0] buf_linear_rsc_dat;
  input buf_linear_rsc_vld;
  output buf_linear_rsc_rdy;
  input core_wen;
  input buf_linear_rsci_oswt_unreg;
  output buf_linear_rsci_bawt;
  input buf_linear_rsci_iswt0;
  output buf_linear_rsci_wen_comp;
  output [4031:0] buf_linear_rsci_idat_mxwt;


  // Interconnect Declarations
  wire buf_linear_rsci_biwt;
  wire buf_linear_rsci_bdwt;
  wire buf_linear_rsci_bcwt;
  wire buf_linear_rsci_irdy_core_sct;
  wire buf_linear_rsci_ivld;
  wire [4031:0] buf_linear_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd16),
  .width(32'sd4032)) buf_linear_rsci (
      .rdy(buf_linear_rsc_rdy),
      .vld(buf_linear_rsc_vld),
      .dat(buf_linear_rsc_dat),
      .irdy(buf_linear_rsci_irdy_core_sct),
      .ivld(buf_linear_rsci_ivld),
      .idat(buf_linear_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci_buf_linear_wait_ctrl
      compute_core_buf_linear_rsci_buf_linear_wait_ctrl_inst (
      .core_wen(core_wen),
      .buf_linear_rsci_oswt_unreg(buf_linear_rsci_oswt_unreg),
      .buf_linear_rsci_iswt0(buf_linear_rsci_iswt0),
      .buf_linear_rsci_biwt(buf_linear_rsci_biwt),
      .buf_linear_rsci_bdwt(buf_linear_rsci_bdwt),
      .buf_linear_rsci_bcwt(buf_linear_rsci_bcwt),
      .buf_linear_rsci_irdy_core_sct(buf_linear_rsci_irdy_core_sct),
      .buf_linear_rsci_ivld(buf_linear_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci_buf_linear_wait_dp compute_core_buf_linear_rsci_buf_linear_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .buf_linear_rsci_oswt_unreg(buf_linear_rsci_oswt_unreg),
      .buf_linear_rsci_bawt(buf_linear_rsci_bawt),
      .buf_linear_rsci_wen_comp(buf_linear_rsci_wen_comp),
      .buf_linear_rsci_idat_mxwt(buf_linear_rsci_idat_mxwt),
      .buf_linear_rsci_biwt(buf_linear_rsci_biwt),
      .buf_linear_rsci_bdwt(buf_linear_rsci_bdwt),
      .buf_linear_rsci_bcwt(buf_linear_rsci_bcwt),
      .buf_linear_rsci_idat(buf_linear_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt_unreg,
      conf_info_rsci_bawt, conf_info_rsci_iswt0, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;
  wire [63:0] conf_info_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd15),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_ctrl compute_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_iswt0(conf_info_rsci_iswt0),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_dp compute_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt_pconst),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
  assign conf_info_rsci_idat_mxwt = conf_info_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt_unreg, done_rsci_bawt,
      done_rsci_iswt0, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  input done_rsci_iswt0;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd27)) done_rsci
      (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci_done_wait_ctrl store_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_iswt0(done_rsci_iswt0),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci_done_wait_dp store_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci (
  clk, rst, dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy,
      core_wen, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_bawt, dma_write_chnl_rsci_iswt0,
      dma_write_chnl_rsci_wen_comp, dma_write_chnl_rsci_idat
);
  input clk;
  input rst;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  input core_wen;
  input dma_write_chnl_rsci_oswt_unreg;
  output dma_write_chnl_rsci_bawt;
  input dma_write_chnl_rsci_iswt0;
  output dma_write_chnl_rsci_wen_comp;
  input [63:0] dma_write_chnl_rsci_idat;


  // Interconnect Declarations
  wire dma_write_chnl_rsci_irdy;
  wire dma_write_chnl_rsci_biwt;
  wire dma_write_chnl_rsci_bdwt;
  wire dma_write_chnl_rsci_bcwt;
  wire dma_write_chnl_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_dma_write_chnl_rsci_idat;
  assign nl_dma_write_chnl_rsci_idat = {32'b11011110101011011011111011101111 , (dma_write_chnl_rsci_idat[31:0])};
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd26),
  .width(32'sd64)) dma_write_chnl_rsci (
      .irdy(dma_write_chnl_rsci_irdy),
      .ivld(dma_write_chnl_rsci_ivld_core_sct),
      .idat(nl_dma_write_chnl_rsci_idat[63:0]),
      .rdy(dma_write_chnl_rsc_rdy),
      .vld(dma_write_chnl_rsc_vld),
      .dat(dma_write_chnl_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
      store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl_inst (
      .core_wen(core_wen),
      .dma_write_chnl_rsci_oswt_unreg(dma_write_chnl_rsci_oswt_unreg),
      .dma_write_chnl_rsci_iswt0(dma_write_chnl_rsci_iswt0),
      .dma_write_chnl_rsci_irdy(dma_write_chnl_rsci_irdy),
      .dma_write_chnl_rsci_biwt(dma_write_chnl_rsci_biwt),
      .dma_write_chnl_rsci_bdwt(dma_write_chnl_rsci_bdwt),
      .dma_write_chnl_rsci_bcwt(dma_write_chnl_rsci_bcwt),
      .dma_write_chnl_rsci_ivld_core_sct(dma_write_chnl_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
      store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_rsci_oswt_unreg(dma_write_chnl_rsci_oswt_unreg),
      .dma_write_chnl_rsci_bawt(dma_write_chnl_rsci_bawt),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .dma_write_chnl_rsci_biwt(dma_write_chnl_rsci_biwt),
      .dma_write_chnl_rsci_bdwt(dma_write_chnl_rsci_bdwt),
      .dma_write_chnl_rsci_bcwt(dma_write_chnl_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci (
  clk, rst, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy,
      core_wen, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_bawt, dma_write_ctrl_rsci_iswt0,
      dma_write_ctrl_rsci_wen_comp, dma_write_ctrl_rsci_idat
);
  input clk;
  input rst;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input core_wen;
  input dma_write_ctrl_rsci_oswt_unreg;
  output dma_write_ctrl_rsci_bawt;
  input dma_write_ctrl_rsci_iswt0;
  output dma_write_ctrl_rsci_wen_comp;
  input [66:0] dma_write_ctrl_rsci_idat;


  // Interconnect Declarations
  wire dma_write_ctrl_rsci_irdy;
  wire dma_write_ctrl_rsci_biwt;
  wire dma_write_ctrl_rsci_bdwt;
  wire dma_write_ctrl_rsci_bcwt;
  wire dma_write_ctrl_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [66:0] nl_dma_write_ctrl_rsci_idat;
  assign nl_dma_write_ctrl_rsci_idat = {51'b011000000000000000000000000000000010000000000000000
      , (dma_write_ctrl_rsci_idat[15:0])};
  esp_acc_conv2dlb_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd25),
  .width(32'sd67)) dma_write_ctrl_rsci (
      .irdy(dma_write_ctrl_rsci_irdy),
      .ivld(dma_write_ctrl_rsci_ivld_core_sct),
      .idat(nl_dma_write_ctrl_rsci_idat[66:0]),
      .rdy(dma_write_ctrl_rsc_rdy),
      .vld(dma_write_ctrl_rsc_vld),
      .dat(dma_write_ctrl_rsc_dat)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
      store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl_inst (
      .core_wen(core_wen),
      .dma_write_ctrl_rsci_oswt_unreg(dma_write_ctrl_rsci_oswt_unreg),
      .dma_write_ctrl_rsci_iswt0(dma_write_ctrl_rsci_iswt0),
      .dma_write_ctrl_rsci_irdy(dma_write_ctrl_rsci_irdy),
      .dma_write_ctrl_rsci_biwt(dma_write_ctrl_rsci_biwt),
      .dma_write_ctrl_rsci_bdwt(dma_write_ctrl_rsci_bdwt),
      .dma_write_ctrl_rsci_bcwt(dma_write_ctrl_rsci_bcwt),
      .dma_write_ctrl_rsci_ivld_core_sct(dma_write_ctrl_rsci_ivld_core_sct)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
      store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_rsci_oswt_unreg(dma_write_ctrl_rsci_oswt_unreg),
      .dma_write_ctrl_rsci_bawt(dma_write_ctrl_rsci_bawt),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_ctrl_rsci_biwt(dma_write_ctrl_rsci_biwt),
      .dma_write_ctrl_rsci_bdwt(dma_write_ctrl_rsci_bdwt),
      .dma_write_ctrl_rsci_bcwt(dma_write_ctrl_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci (
  clk, rst, var_output_rsc_dat, var_output_rsc_vld, var_output_rsc_rdy, core_wen,
      var_output_rsci_oswt_unreg, var_output_rsci_bawt, var_output_rsci_iswt0, var_output_rsci_wen_comp,
      var_output_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [31:0] var_output_rsc_dat;
  input var_output_rsc_vld;
  output var_output_rsc_rdy;
  input core_wen;
  input var_output_rsci_oswt_unreg;
  output var_output_rsci_bawt;
  input var_output_rsci_iswt0;
  output var_output_rsci_wen_comp;
  output [31:0] var_output_rsci_idat_mxwt;


  // Interconnect Declarations
  wire var_output_rsci_biwt;
  wire var_output_rsci_bdwt;
  wire var_output_rsci_bcwt;
  wire var_output_rsci_irdy_core_sct;
  wire var_output_rsci_ivld;
  wire [31:0] var_output_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd24),
  .width(32'sd32)) var_output_rsci (
      .rdy(var_output_rsc_rdy),
      .vld(var_output_rsc_vld),
      .dat(var_output_rsc_dat),
      .irdy(var_output_rsci_irdy_core_sct),
      .ivld(var_output_rsci_ivld),
      .idat(var_output_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci_var_output_wait_ctrl store_core_var_output_rsci_var_output_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .var_output_rsci_oswt_unreg(var_output_rsci_oswt_unreg),
      .var_output_rsci_iswt0(var_output_rsci_iswt0),
      .var_output_rsci_biwt(var_output_rsci_biwt),
      .var_output_rsci_bdwt(var_output_rsci_bdwt),
      .var_output_rsci_bcwt(var_output_rsci_bcwt),
      .var_output_rsci_irdy_core_sct(var_output_rsci_irdy_core_sct),
      .var_output_rsci_ivld(var_output_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci_var_output_wait_dp store_core_var_output_rsci_var_output_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .var_output_rsci_oswt_unreg(var_output_rsci_oswt_unreg),
      .var_output_rsci_bawt(var_output_rsci_bawt),
      .var_output_rsci_wen_comp(var_output_rsci_wen_comp),
      .var_output_rsci_idat_mxwt(var_output_rsci_idat_mxwt),
      .var_output_rsci_biwt(var_output_rsci_biwt),
      .var_output_rsci_bdwt(var_output_rsci_bdwt),
      .var_output_rsci_bcwt(var_output_rsci_bcwt),
      .var_output_rsci_idat(var_output_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt_unreg,
      conf_info_rsci_bawt, conf_info_rsci_iswt0, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;
  wire [63:0] conf_info_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd23),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_ctrl store_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_iswt0(conf_info_rsci_iswt0),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_dp store_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt_pconst),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
  assign conf_info_rsci_idat_mxwt = conf_info_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core (
  clk, rst, acc_done_rsc_vld, config_done_cns_rdy, config_done_cns_vld, load_done_cns_rdy,
      load_done_cns_vld, compute_done_cns_rdy, compute_done_cns_vld, store_done_cns_rdy,
      store_done_cns_vld
);
  input clk;
  input rst;
  output acc_done_rsc_vld;
  output config_done_cns_rdy;
  input config_done_cns_vld;
  output load_done_cns_rdy;
  input load_done_cns_vld;
  output compute_done_cns_rdy;
  input compute_done_cns_vld;
  output store_done_cns_rdy;
  input store_done_cns_vld;


  // Interconnect Declarations
  wire core_wen;
  wire acc_done_rsci_bawt;
  wire core_wten;
  wire config_done_cnsi_bawt;
  wire config_done_cnsi_wen_comp;
  wire load_done_cnsi_bawt;
  wire load_done_cnsi_wen_comp;
  reg load_done_cnsi_irdy_core_psct;
  wire compute_done_cnsi_bawt;
  wire compute_done_cnsi_wen_comp;
  wire store_done_cnsi_bawt;
  wire store_done_cnsi_wen_comp;
  wire [1:0] fsm_output;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_5;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_21;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_56_cse;
  reg main_stage_v_4;
  reg reg_store_done_cnsi_irdy_core_psct_cse;
  reg reg_compute_done_cnsi_irdy_core_psct_cse;
  reg reg_store_done_cnsi_oswt_cse;
  reg reg_load_done_cnsi_iswt0_cse;
  wire or_20_cse;
  wire or_17_cse;
  wire or_15_cse;
  wire or_cse;
  wire main_stage_v_4_mx0c1;
  reg reg_config_done_cnsi_iswt0_cse;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_acc_done_rsci conv2dlb_cxx_catapult_core_core_acc_done_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .acc_done_rsc_vld(acc_done_rsc_vld),
      .core_wen(core_wen),
      .acc_done_rsci_oswt_unreg(and_dcpl_27),
      .acc_done_rsci_bawt(acc_done_rsci_bawt),
      .acc_done_rsci_iswt0(reg_store_done_cnsi_oswt_cse),
      .core_wten(core_wten)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_config_done_cnsi
      conv2dlb_cxx_catapult_core_core_config_done_cnsi_inst (
      .clk(clk),
      .rst(rst),
      .config_done_cns_rdy(config_done_cns_rdy),
      .config_done_cns_vld(config_done_cns_vld),
      .core_wen(core_wen),
      .config_done_cnsi_oswt_unreg(and_56_cse),
      .config_done_cnsi_bawt(config_done_cnsi_bawt),
      .config_done_cnsi_iswt0(reg_config_done_cnsi_iswt0_cse),
      .config_done_cnsi_wen_comp(config_done_cnsi_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_load_done_cnsi conv2dlb_cxx_catapult_core_core_load_done_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .load_done_cns_rdy(load_done_cns_rdy),
      .load_done_cns_vld(load_done_cns_vld),
      .core_wen(core_wen),
      .load_done_cnsi_oswt_unreg(and_dcpl_19),
      .load_done_cnsi_bawt(load_done_cnsi_bawt),
      .load_done_cnsi_iswt0(reg_load_done_cnsi_iswt0_cse),
      .load_done_cnsi_wen_comp(load_done_cnsi_wen_comp),
      .load_done_cnsi_irdy_core_psct(load_done_cnsi_irdy_core_psct)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_compute_done_cnsi
      conv2dlb_cxx_catapult_core_core_compute_done_cnsi_inst (
      .clk(clk),
      .rst(rst),
      .compute_done_cns_rdy(compute_done_cns_rdy),
      .compute_done_cns_vld(compute_done_cns_vld),
      .core_wen(core_wen),
      .compute_done_cnsi_oswt_unreg(and_dcpl_14),
      .compute_done_cnsi_bawt(compute_done_cnsi_bawt),
      .compute_done_cnsi_iswt0(reg_compute_done_cnsi_irdy_core_psct_cse),
      .compute_done_cnsi_wen_comp(compute_done_cnsi_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_store_done_cnsi conv2dlb_cxx_catapult_core_core_store_done_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .store_done_cns_rdy(store_done_cns_rdy),
      .store_done_cns_vld(store_done_cns_vld),
      .core_wen(core_wen),
      .store_done_cnsi_oswt_unreg(and_dcpl_18),
      .store_done_cnsi_bawt(store_done_cnsi_bawt),
      .store_done_cnsi_iswt0(reg_store_done_cnsi_irdy_core_psct_cse),
      .store_done_cnsi_wen_comp(store_done_cnsi_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_staller conv2dlb_cxx_catapult_core_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .config_done_cnsi_wen_comp(config_done_cnsi_wen_comp),
      .load_done_cnsi_wen_comp(load_done_cnsi_wen_comp),
      .compute_done_cnsi_wen_comp(compute_done_cnsi_wen_comp),
      .store_done_cnsi_wen_comp(store_done_cnsi_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core_core_fsm conv2dlb_cxx_catapult_core_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_20_cse = load_done_cnsi_bawt | (~ reg_load_done_cnsi_iswt0_cse);
  assign or_17_cse = compute_done_cnsi_bawt | (~ reg_compute_done_cnsi_irdy_core_psct_cse);
  assign or_15_cse = store_done_cnsi_bawt | (~ reg_store_done_cnsi_irdy_core_psct_cse);
  assign or_cse = acc_done_rsci_bawt | (~ main_stage_v_4);
  assign and_dcpl_1 = or_cse & or_15_cse;
  assign and_dcpl_2 = and_dcpl_1 & or_17_cse;
  assign and_dcpl_5 = load_done_cnsi_bawt & reg_load_done_cnsi_iswt0_cse;
  assign and_dcpl_13 = compute_done_cnsi_bawt & reg_compute_done_cnsi_irdy_core_psct_cse;
  assign and_dcpl_14 = and_dcpl_1 & and_dcpl_13;
  assign and_dcpl_17 = or_cse & store_done_cnsi_bawt & (~(compute_done_cnsi_bawt
      & reg_compute_done_cnsi_irdy_core_psct_cse)) & reg_store_done_cnsi_irdy_core_psct_cse;
  assign and_dcpl_18 = or_cse & reg_store_done_cnsi_irdy_core_psct_cse & store_done_cnsi_bawt;
  assign and_dcpl_19 = and_dcpl_2 & and_dcpl_5;
  assign and_dcpl_21 = and_dcpl_1 & and_dcpl_13 & (~(load_done_cnsi_bawt & reg_load_done_cnsi_iswt0_cse));
  assign and_dcpl_26 = and_dcpl_2 & and_dcpl_5 & (~ config_done_cnsi_bawt);
  assign and_dcpl_27 = main_stage_v_4 & acc_done_rsci_bawt;
  assign and_56_cse = and_dcpl_2 & or_20_cse & config_done_cnsi_bawt & (fsm_output[1]);
  assign main_stage_v_4_mx0c1 = and_dcpl_27 & (~(store_done_cnsi_bawt & reg_store_done_cnsi_irdy_core_psct_cse));
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_config_done_cnsi_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((config_done_cnsi_bawt & or_20_cse & or_17_cse & or_15_cse
        & or_cse) | (fsm_output[0])) ) begin
      reg_config_done_cnsi_iswt0_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_store_done_cnsi_irdy_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_14 | and_dcpl_17) ) begin
      reg_store_done_cnsi_irdy_core_psct_cse <= ~ and_dcpl_17;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_store_done_cnsi_oswt_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_store_done_cnsi_oswt_cse <= and_dcpl_18;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_compute_done_cnsi_irdy_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_19 | and_dcpl_21) ) begin
      reg_compute_done_cnsi_irdy_core_psct_cse <= ~ and_dcpl_21;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      load_done_cnsi_irdy_core_psct <= 1'b0;
    end
    else if ( core_wen & (and_56_cse | (and_dcpl_2 & and_dcpl_5 & config_done_cnsi_bawt)
        | and_dcpl_26) ) begin
      load_done_cnsi_irdy_core_psct <= ~ and_dcpl_26;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_load_done_cnsi_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (and_56_cse | and_dcpl_26) ) begin
      reg_load_done_cnsi_iswt0_cse <= ~ and_dcpl_26;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_18 | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config_core
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_conf_load_rsc_dat,
      plm_conf_load_rsc_vld, plm_conf_load_rsc_rdy, plm_conf_compute_rsc_dat, plm_conf_compute_rsc_vld,
      plm_conf_compute_rsc_rdy, plm_conf_store_rsc_dat, plm_conf_store_rsc_vld, plm_conf_store_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [255:0] plm_conf_load_rsc_dat;
  output plm_conf_load_rsc_vld;
  input plm_conf_load_rsc_rdy;
  output [255:0] plm_conf_compute_rsc_dat;
  output plm_conf_compute_rsc_vld;
  input plm_conf_compute_rsc_rdy;
  output [255:0] plm_conf_store_rsc_dat;
  output plm_conf_store_rsc_vld;
  input plm_conf_store_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire core_wen;
  wire conf_info_rsci_bawt;
  wire conf_info_rsci_wen_comp;
  wire [255:0] conf_info_rsci_idat_mxwt;
  wire plm_conf_load_rsci_bawt;
  wire plm_conf_load_rsci_wen_comp;
  wire plm_conf_compute_rsci_bawt;
  wire plm_conf_compute_rsci_wen_comp;
  wire plm_conf_store_rsci_bawt;
  wire plm_conf_store_rsci_wen_comp;
  reg [255:0] plm_conf_store_rsci_idat;
  wire done_rsci_bawt;
  wire done_rsci_wen_comp;
  wire [1:0] fsm_output;
  wire and_dcpl_1;
  wire and_dcpl_9;
  wire or_dcpl_3;
  wire or_dcpl_5;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire or_dcpl_6;
  wire and_dcpl_17;
  wire and_dcpl_20;
  wire or_tmp_8;
  reg reg_done_rsci_ivld_core_psct_cse;
  reg reg_plm_conf_store_rsci_ivld_core_psct_cse;
  reg [255:0] reg_plm_conf_compute_rsci_idat_cse;
  wire or_cse;
  reg reg_conf_info_rsci_iswt0_cse;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_config_core_conf_info_rsci config_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(or_tmp_8),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_iswt0(reg_conf_info_rsci_iswt0_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_load_rsci config_core_plm_conf_load_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_conf_load_rsc_dat(plm_conf_load_rsc_dat),
      .plm_conf_load_rsc_vld(plm_conf_load_rsc_vld),
      .plm_conf_load_rsc_rdy(plm_conf_load_rsc_rdy),
      .core_wen(core_wen),
      .plm_conf_load_rsci_oswt_unreg(and_dcpl_15),
      .plm_conf_load_rsci_bawt(plm_conf_load_rsci_bawt),
      .plm_conf_load_rsci_iswt0(reg_plm_conf_store_rsci_ivld_core_psct_cse),
      .plm_conf_load_rsci_wen_comp(plm_conf_load_rsci_wen_comp),
      .plm_conf_load_rsci_idat(reg_plm_conf_compute_rsci_idat_cse)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_compute_rsci config_core_plm_conf_compute_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_conf_compute_rsc_dat(plm_conf_compute_rsc_dat),
      .plm_conf_compute_rsc_vld(plm_conf_compute_rsc_vld),
      .plm_conf_compute_rsc_rdy(plm_conf_compute_rsc_rdy),
      .core_wen(core_wen),
      .plm_conf_compute_rsci_oswt_unreg(and_dcpl_15),
      .plm_conf_compute_rsci_bawt(plm_conf_compute_rsci_bawt),
      .plm_conf_compute_rsci_iswt0(reg_plm_conf_store_rsci_ivld_core_psct_cse),
      .plm_conf_compute_rsci_wen_comp(plm_conf_compute_rsci_wen_comp),
      .plm_conf_compute_rsci_idat(reg_plm_conf_compute_rsci_idat_cse)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_plm_conf_store_rsci config_core_plm_conf_store_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_conf_store_rsc_dat(plm_conf_store_rsc_dat),
      .plm_conf_store_rsc_vld(plm_conf_store_rsc_vld),
      .plm_conf_store_rsc_rdy(plm_conf_store_rsc_rdy),
      .core_wen(core_wen),
      .plm_conf_store_rsci_oswt_unreg(and_dcpl_15),
      .plm_conf_store_rsci_bawt(plm_conf_store_rsci_bawt),
      .plm_conf_store_rsci_iswt0(reg_plm_conf_store_rsci_ivld_core_psct_cse),
      .plm_conf_store_rsci_wen_comp(plm_conf_store_rsci_wen_comp),
      .plm_conf_store_rsci_idat(plm_conf_store_rsci_idat)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_done_rsci config_core_done_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(and_dcpl_16),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_iswt0(reg_done_rsci_ivld_core_psct_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_staller config_core_staller_inst (
      .core_wen(core_wen),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .plm_conf_load_rsci_wen_comp(plm_conf_load_rsci_wen_comp),
      .plm_conf_compute_rsci_wen_comp(plm_conf_compute_rsci_wen_comp),
      .plm_conf_store_rsci_wen_comp(plm_conf_store_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_config_core_core_fsm config_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_cse = done_rsci_bawt | (~ reg_done_rsci_ivld_core_psct_cse);
  assign and_dcpl_1 = plm_conf_load_rsci_bawt & plm_conf_compute_rsci_bawt;
  assign and_dcpl_9 = reg_done_rsci_ivld_core_psct_cse & (~ done_rsci_bawt);
  assign or_dcpl_3 = ~(plm_conf_load_rsci_bawt & plm_conf_compute_rsci_bawt);
  assign or_dcpl_5 = ((or_dcpl_3 | (~ plm_conf_store_rsci_bawt)) & reg_plm_conf_store_rsci_ivld_core_psct_cse)
      | and_dcpl_9 | (~ conf_info_rsci_bawt);
  assign and_dcpl_15 = or_cse & plm_conf_load_rsci_bawt & plm_conf_compute_rsci_bawt
      & plm_conf_store_rsci_bawt & reg_plm_conf_store_rsci_ivld_core_psct_cse;
  assign and_dcpl_16 = reg_done_rsci_ivld_core_psct_cse & done_rsci_bawt;
  assign or_dcpl_6 = ~(plm_conf_store_rsci_bawt & reg_plm_conf_store_rsci_ivld_core_psct_cse);
  assign and_dcpl_17 = (or_dcpl_3 | or_dcpl_6) & and_dcpl_16;
  assign and_dcpl_20 = or_cse & and_dcpl_1 & plm_conf_store_rsci_bawt & reg_plm_conf_store_rsci_ivld_core_psct_cse
      & (~ conf_info_rsci_bawt);
  assign or_tmp_8 = (~((~(and_dcpl_1 & plm_conf_store_rsci_bawt)) & reg_plm_conf_store_rsci_ivld_core_psct_cse))
      & or_cse & conf_info_rsci_bawt & (fsm_output[1]);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((conf_info_rsci_bawt & (plm_conf_load_rsci_bawt | (~ reg_plm_conf_store_rsci_ivld_core_psct_cse))
        & (plm_conf_compute_rsci_bawt | (~ reg_plm_conf_store_rsci_ivld_core_psct_cse))
        & (plm_conf_store_rsci_bawt | (~ reg_plm_conf_store_rsci_ivld_core_psct_cse))
        & or_cse) | (fsm_output[0])) ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_done_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_15 | and_dcpl_17) ) begin
      reg_done_rsci_ivld_core_psct_cse <= ~ and_dcpl_17;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_store_rsci_idat <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_5 | ((and_dcpl_9 | or_dcpl_3 | or_dcpl_6 | (~
        conf_info_rsci_bawt)) & (fsm_output[0])))) ) begin
      plm_conf_store_rsci_idat <= conf_info_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_conf_store_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_8 | and_dcpl_20) ) begin
      reg_plm_conf_store_rsci_ivld_core_psct_cse <= ~ and_dcpl_20;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_conf_compute_rsci_idat_cse <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_5 | (fsm_output[0]))) ) begin
      reg_plm_conf_compute_rsci_idat_cse <= conf_info_rsci_idat_mxwt;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load_core
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, buf_linear_rsc_dat,
      buf_linear_rsc_vld, buf_linear_rsc_rdy, plm_kernel_rsc_dat, plm_kernel_rsc_vld,
      plm_kernel_rsc_rdy, dma_read_ctrl_rsc_dat, dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy,
      dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy, done_rsc_rdy,
      done_rsc_vld, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d, LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [4031:0] buf_linear_rsc_dat;
  output buf_linear_rsc_vld;
  input buf_linear_rsc_rdy;
  output [1567:0] plm_kernel_rsc_dat;
  output plm_kernel_rsc_vld;
  input plm_kernel_rsc_rdy;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;
  output [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d;
  input [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d;
  output [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d;
  output [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire conf_info_rsci_wen_comp;
  wire [231:0] conf_info_rsci_idat_mxwt;
  wire buf_linear_rsci_bawt;
  wire buf_linear_rsci_wen_comp;
  wire plm_kernel_rsci_bawt;
  wire plm_kernel_rsci_wen_comp;
  wire dma_read_ctrl_rsci_bawt;
  wire dma_read_ctrl_rsci_irdy_mxwt;
  wire dma_read_chnl_rsci_bawt;
  wire dma_read_chnl_rsci_wen_comp;
  wire [31:0] dma_read_chnl_rsci_idat_mxwt;
  wire done_rsci_wen_comp;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt;
  wire [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt;
  reg [31:0] buf_linear_rsci_idat_4031_4000;
  reg [31:0] buf_linear_rsci_idat_3999_3968;
  reg [31:0] buf_linear_rsci_idat_3967_3936;
  reg [31:0] buf_linear_rsci_idat_3935_3904;
  reg [31:0] buf_linear_rsci_idat_3903_3872;
  reg [31:0] buf_linear_rsci_idat_3871_3840;
  reg [31:0] buf_linear_rsci_idat_3839_3808;
  reg [31:0] buf_linear_rsci_idat_3807_3776;
  reg [31:0] buf_linear_rsci_idat_3775_3744;
  reg [31:0] buf_linear_rsci_idat_3743_3712;
  reg [31:0] buf_linear_rsci_idat_3711_3680;
  reg [31:0] buf_linear_rsci_idat_3679_3648;
  reg [31:0] buf_linear_rsci_idat_3647_3616;
  reg [31:0] buf_linear_rsci_idat_3615_3584;
  reg [31:0] buf_linear_rsci_idat_3583_3552;
  reg [31:0] buf_linear_rsci_idat_3551_3520;
  reg [31:0] buf_linear_rsci_idat_3519_3488;
  reg [31:0] buf_linear_rsci_idat_3487_3456;
  reg [31:0] buf_linear_rsci_idat_3455_3424;
  reg [31:0] buf_linear_rsci_idat_3423_3392;
  reg [31:0] buf_linear_rsci_idat_3391_3360;
  reg [31:0] buf_linear_rsci_idat_3359_3328;
  reg [31:0] buf_linear_rsci_idat_3327_3296;
  reg [31:0] buf_linear_rsci_idat_3295_3264;
  reg [31:0] buf_linear_rsci_idat_3263_3232;
  reg [31:0] buf_linear_rsci_idat_3231_3200;
  reg [31:0] buf_linear_rsci_idat_3199_3168;
  reg [31:0] buf_linear_rsci_idat_3167_3136;
  reg [31:0] buf_linear_rsci_idat_3135_3104;
  reg [31:0] buf_linear_rsci_idat_3103_3072;
  reg [31:0] buf_linear_rsci_idat_3071_3040;
  reg [31:0] buf_linear_rsci_idat_3039_3008;
  reg [31:0] buf_linear_rsci_idat_3007_2976;
  reg [31:0] buf_linear_rsci_idat_2975_2944;
  reg [31:0] buf_linear_rsci_idat_2943_2912;
  reg [31:0] buf_linear_rsci_idat_2911_2880;
  reg [31:0] buf_linear_rsci_idat_2879_2848;
  reg [31:0] buf_linear_rsci_idat_2847_2816;
  reg [31:0] buf_linear_rsci_idat_2815_2784;
  reg [31:0] buf_linear_rsci_idat_2783_2752;
  reg [31:0] buf_linear_rsci_idat_2751_2720;
  reg [31:0] buf_linear_rsci_idat_2719_2688;
  reg [31:0] buf_linear_rsci_idat_2687_2656;
  reg [31:0] buf_linear_rsci_idat_2655_2624;
  reg [31:0] buf_linear_rsci_idat_2623_2592;
  reg [31:0] buf_linear_rsci_idat_2591_2560;
  reg [31:0] buf_linear_rsci_idat_2559_2528;
  reg [31:0] buf_linear_rsci_idat_2527_2496;
  reg [31:0] buf_linear_rsci_idat_2495_2464;
  reg [31:0] buf_linear_rsci_idat_2463_2432;
  reg [31:0] buf_linear_rsci_idat_2431_2400;
  reg [31:0] buf_linear_rsci_idat_2399_2368;
  reg [31:0] buf_linear_rsci_idat_2367_2336;
  reg [31:0] buf_linear_rsci_idat_2335_2304;
  reg [31:0] buf_linear_rsci_idat_2303_2272;
  reg [31:0] buf_linear_rsci_idat_2271_2240;
  reg [31:0] buf_linear_rsci_idat_2239_2208;
  reg [31:0] buf_linear_rsci_idat_2207_2176;
  reg [31:0] buf_linear_rsci_idat_2175_2144;
  reg [31:0] buf_linear_rsci_idat_2143_2112;
  reg [31:0] buf_linear_rsci_idat_2111_2080;
  reg [31:0] buf_linear_rsci_idat_2079_2048;
  reg [31:0] buf_linear_rsci_idat_2047_2016;
  reg [31:0] buf_linear_rsci_idat_2015_1984;
  reg [31:0] buf_linear_rsci_idat_1983_1952;
  reg [31:0] buf_linear_rsci_idat_1951_1920;
  reg [31:0] buf_linear_rsci_idat_1919_1888;
  reg [31:0] buf_linear_rsci_idat_1887_1856;
  reg [31:0] buf_linear_rsci_idat_1855_1824;
  reg [31:0] buf_linear_rsci_idat_1823_1792;
  reg [31:0] buf_linear_rsci_idat_1791_1760;
  reg [31:0] buf_linear_rsci_idat_1759_1728;
  reg [31:0] buf_linear_rsci_idat_1727_1696;
  reg [31:0] buf_linear_rsci_idat_1695_1664;
  reg [31:0] buf_linear_rsci_idat_1663_1632;
  reg [31:0] buf_linear_rsci_idat_1631_1600;
  reg [31:0] buf_linear_rsci_idat_1599_1568;
  reg [31:0] buf_linear_rsci_idat_1567_1536;
  reg [31:0] buf_linear_rsci_idat_1535_1504;
  reg [31:0] buf_linear_rsci_idat_1503_1472;
  reg [31:0] buf_linear_rsci_idat_1471_1440;
  reg [31:0] buf_linear_rsci_idat_1439_1408;
  reg [31:0] buf_linear_rsci_idat_1407_1376;
  reg [31:0] buf_linear_rsci_idat_1375_1344;
  reg [31:0] buf_linear_rsci_idat_1343_1312;
  reg [31:0] buf_linear_rsci_idat_1311_1280;
  reg [31:0] buf_linear_rsci_idat_1279_1248;
  reg [31:0] buf_linear_rsci_idat_1247_1216;
  reg [31:0] buf_linear_rsci_idat_1215_1184;
  reg [31:0] buf_linear_rsci_idat_1183_1152;
  reg [31:0] buf_linear_rsci_idat_1151_1120;
  reg [31:0] buf_linear_rsci_idat_1119_1088;
  reg [31:0] buf_linear_rsci_idat_1087_1056;
  reg [31:0] buf_linear_rsci_idat_1055_1024;
  reg [31:0] buf_linear_rsci_idat_1023_992;
  reg [31:0] buf_linear_rsci_idat_991_960;
  reg [31:0] buf_linear_rsci_idat_959_928;
  reg [31:0] buf_linear_rsci_idat_927_896;
  reg [31:0] buf_linear_rsci_idat_895_864;
  reg [31:0] buf_linear_rsci_idat_863_832;
  reg [31:0] buf_linear_rsci_idat_831_800;
  reg [31:0] buf_linear_rsci_idat_799_768;
  reg [31:0] buf_linear_rsci_idat_767_736;
  reg [31:0] buf_linear_rsci_idat_735_704;
  reg [31:0] buf_linear_rsci_idat_703_672;
  reg [31:0] buf_linear_rsci_idat_671_640;
  reg [31:0] buf_linear_rsci_idat_639_608;
  reg [31:0] buf_linear_rsci_idat_607_576;
  reg [31:0] buf_linear_rsci_idat_575_544;
  reg [31:0] buf_linear_rsci_idat_543_512;
  reg [31:0] buf_linear_rsci_idat_511_480;
  reg [31:0] buf_linear_rsci_idat_479_448;
  reg [31:0] buf_linear_rsci_idat_447_416;
  reg [31:0] buf_linear_rsci_idat_415_384;
  reg [31:0] buf_linear_rsci_idat_383_352;
  reg [31:0] buf_linear_rsci_idat_351_320;
  reg [31:0] buf_linear_rsci_idat_319_288;
  reg [31:0] buf_linear_rsci_idat_287_256;
  reg [31:0] buf_linear_rsci_idat_255_224;
  reg [31:0] buf_linear_rsci_idat_223_192;
  reg [31:0] buf_linear_rsci_idat_191_160;
  reg [31:0] buf_linear_rsci_idat_159_128;
  reg [31:0] buf_linear_rsci_idat_127_96;
  reg [31:0] buf_linear_rsci_idat_95_64;
  reg [31:0] buf_linear_rsci_idat_63_32;
  reg [31:0] buf_linear_rsci_idat_31_0;
  reg [31:0] plm_kernel_rsci_idat_1567_1536;
  reg [31:0] plm_kernel_rsci_idat_1535_1504;
  reg [31:0] plm_kernel_rsci_idat_1503_1472;
  reg [31:0] plm_kernel_rsci_idat_1471_1440;
  reg [31:0] plm_kernel_rsci_idat_1439_1408;
  reg [31:0] plm_kernel_rsci_idat_1407_1376;
  reg [31:0] plm_kernel_rsci_idat_1375_1344;
  reg [31:0] plm_kernel_rsci_idat_1343_1312;
  reg [31:0] plm_kernel_rsci_idat_1311_1280;
  reg [31:0] plm_kernel_rsci_idat_1279_1248;
  reg [31:0] plm_kernel_rsci_idat_1247_1216;
  reg [31:0] plm_kernel_rsci_idat_1215_1184;
  reg [31:0] plm_kernel_rsci_idat_1183_1152;
  reg [31:0] plm_kernel_rsci_idat_1151_1120;
  reg [31:0] plm_kernel_rsci_idat_1119_1088;
  reg [31:0] plm_kernel_rsci_idat_1087_1056;
  reg [31:0] plm_kernel_rsci_idat_1055_1024;
  reg [31:0] plm_kernel_rsci_idat_1023_992;
  reg [31:0] plm_kernel_rsci_idat_991_960;
  reg [31:0] plm_kernel_rsci_idat_959_928;
  reg [31:0] plm_kernel_rsci_idat_927_896;
  reg [31:0] plm_kernel_rsci_idat_895_864;
  reg [31:0] plm_kernel_rsci_idat_863_832;
  reg [31:0] plm_kernel_rsci_idat_831_800;
  reg [31:0] plm_kernel_rsci_idat_799_768;
  reg [31:0] plm_kernel_rsci_idat_767_736;
  reg [31:0] plm_kernel_rsci_idat_735_704;
  reg [31:0] plm_kernel_rsci_idat_703_672;
  reg [31:0] plm_kernel_rsci_idat_671_640;
  reg [31:0] plm_kernel_rsci_idat_639_608;
  reg [31:0] plm_kernel_rsci_idat_607_576;
  reg [31:0] plm_kernel_rsci_idat_575_544;
  reg [31:0] plm_kernel_rsci_idat_543_512;
  reg [31:0] plm_kernel_rsci_idat_511_480;
  reg [31:0] plm_kernel_rsci_idat_479_448;
  reg [31:0] plm_kernel_rsci_idat_447_416;
  reg [31:0] plm_kernel_rsci_idat_415_384;
  reg [31:0] plm_kernel_rsci_idat_383_352;
  reg [31:0] plm_kernel_rsci_idat_351_320;
  reg [31:0] plm_kernel_rsci_idat_319_288;
  reg [31:0] plm_kernel_rsci_idat_287_256;
  reg [31:0] plm_kernel_rsci_idat_255_224;
  reg [31:0] plm_kernel_rsci_idat_223_192;
  reg [31:0] plm_kernel_rsci_idat_191_160;
  reg [31:0] plm_kernel_rsci_idat_159_128;
  reg [31:0] plm_kernel_rsci_idat_127_96;
  reg [31:0] plm_kernel_rsci_idat_95_64;
  reg [31:0] plm_kernel_rsci_idat_63_32;
  reg [31:0] plm_kernel_rsci_idat_31_0;
  reg [15:0] dma_read_ctrl_rsci_idat_47_32;
  reg [15:0] dma_read_ctrl_rsci_idat_15_0;
  wire [3:0] fsm_output;
  wire [4:0] LOAD_BATCH_LOOP_acc_tmp;
  wire [5:0] nl_LOAD_BATCH_LOOP_acc_tmp;
  wire LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_nor_tmp;
  wire [5:0] LOAD_LOOP_acc_tmp;
  wire [6:0] nl_LOAD_LOOP_acc_tmp;
  wire LOAD_LOOP_if_equal_tmp;
  wire [8:0] operator_8_false_7_acc_tmp;
  wire [9:0] nl_operator_8_false_7_acc_tmp;
  wire LOAD_LOOP_for_if_for_for_if_equal_tmp;
  wire [8:0] operator_8_false_1_acc_tmp;
  wire [9:0] nl_operator_8_false_1_acc_tmp;
  wire [5:0] LOAD_LOOP_for_acc_2_tmp;
  wire [6:0] nl_LOAD_LOOP_for_acc_2_tmp;
  wire LOAD_LOOP_for_if_3_equal_tmp;
  wire [8:0] operator_8_false_6_acc_tmp;
  wire [9:0] nl_operator_8_false_6_acc_tmp;
  wire LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_1_LOAD_LOOP_for_if_2_for_if_1_nor_tmp;
  wire LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_if_1_LOAD_LOOP_for_if_2_for_for_if_1_nor_tmp;
  wire LOAD_BATCH_LOOP_and_4_tmp;
  wire [1:0] LOAD_LOOP_for_if_2_for_mux1h_378_tmp;
  wire LOAD_BATCH_LOOP_and_3_tmp;
  wire or_tmp_4;
  wire or_tmp_57;
  wire and_tmp_12;
  wire or_tmp_90;
  wire mux_tmp_52;
  wire nor_tmp_50;
  wire mux_tmp_80;
  wire and_dcpl_24;
  wire nor_tmp_54;
  wire or_tmp_148;
  wire and_tmp_17;
  wire or_tmp_151;
  wire mux_tmp_91;
  wire mux_tmp_93;
  wire and_dcpl_28;
  wire or_tmp_154;
  wire mux_tmp_103;
  wire nor_tmp_63;
  wire mux_tmp_109;
  wire nor_tmp_67;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire and_dcpl_44;
  wire or_dcpl_29;
  wire or_dcpl_30;
  wire or_dcpl_31;
  wire or_dcpl_32;
  wire or_dcpl_34;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire or_dcpl_38;
  wire or_dcpl_39;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire or_dcpl_41;
  wire or_dcpl_42;
  wire and_dcpl_54;
  wire or_dcpl_44;
  wire or_dcpl_45;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire or_dcpl_47;
  wire and_dcpl_61;
  wire and_dcpl_62;
  wire or_dcpl_49;
  wire and_dcpl_65;
  wire or_dcpl_51;
  wire and_dcpl_68;
  wire or_dcpl_53;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire or_dcpl_55;
  wire or_dcpl_56;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire or_dcpl_65;
  wire or_dcpl_66;
  wire and_dcpl_108;
  wire or_dcpl_76;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire or_dcpl_85;
  wire and_dcpl_144;
  wire or_dcpl_94;
  wire or_dcpl_103;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_172;
  wire and_dcpl_173;
  wire and_dcpl_174;
  wire and_dcpl_176;
  wire and_dcpl_178;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire not_tmp_118;
  wire and_dcpl_186;
  wire and_dcpl_188;
  wire not_tmp_124;
  wire and_dcpl_194;
  wire not_tmp_125;
  wire and_dcpl_200;
  wire not_tmp_126;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_223;
  wire and_dcpl_224;
  wire and_dcpl_241;
  wire and_dcpl_242;
  wire and_dcpl_259;
  wire and_dcpl_260;
  wire and_dcpl_277;
  wire and_dcpl_294;
  wire and_dcpl_311;
  wire and_dcpl_328;
  wire and_dcpl_329;
  wire and_dcpl_330;
  wire and_dcpl_347;
  wire and_dcpl_364;
  wire and_dcpl_381;
  wire and_dcpl_398;
  wire and_dcpl_399;
  wire and_dcpl_416;
  wire and_dcpl_433;
  wire and_dcpl_450;
  wire and_dcpl_467;
  wire and_dcpl_468;
  wire and_dcpl_469;
  wire not_tmp_127;
  wire not_tmp_128;
  wire not_tmp_129;
  wire not_tmp_130;
  wire and_dcpl_486;
  wire and_dcpl_503;
  wire and_dcpl_520;
  wire and_dcpl_537;
  wire and_dcpl_538;
  wire and_dcpl_555;
  wire and_dcpl_572;
  wire and_dcpl_589;
  wire and_dcpl_606;
  wire and_dcpl_607;
  wire and_dcpl_608;
  wire not_tmp_131;
  wire not_tmp_132;
  wire not_tmp_133;
  wire not_tmp_134;
  wire and_dcpl_625;
  wire and_dcpl_642;
  wire and_dcpl_659;
  wire and_dcpl_676;
  wire and_dcpl_677;
  wire not_tmp_135;
  wire not_tmp_136;
  wire not_tmp_137;
  wire not_tmp_138;
  wire and_dcpl_694;
  wire and_dcpl_711;
  wire and_dcpl_728;
  wire and_dcpl_738;
  wire and_dcpl_739;
  wire and_dcpl_752;
  wire or_tmp_325;
  wire nor_tmp_101;
  wire mux_tmp_260;
  wire nand_tmp_29;
  wire or_tmp_340;
  wire and_tmp_22;
  wire nand_tmp_32;
  wire mux_tmp_284;
  wire nand_tmp_34;
  wire or_tmp_352;
  wire and_dcpl_764;
  wire and_dcpl_772;
  wire or_dcpl_122;
  wire or_dcpl_128;
  wire or_dcpl_129;
  wire or_tmp_388;
  wire and_tmp_25;
  wire or_dcpl_135;
  wire or_dcpl_136;
  wire and_dcpl_778;
  wire or_dcpl_146;
  wire and_dcpl_779;
  wire or_tmp_408;
  wire or_tmp_409;
  wire mux_tmp_336;
  wire mux_tmp_338;
  wire mux_tmp_340;
  wire or_dcpl_147;
  wire or_dcpl_150;
  wire mux_tmp_345;
  wire or_tmp_419;
  wire mux_tmp_347;
  wire mux_tmp_349;
  wire mux_tmp_353;
  wire mux_tmp_359;
  wire nand_tmp_41;
  wire or_tmp_471;
  wire and_tmp_30;
  wire and_tmp_32;
  wire nor_tmp_172;
  wire nor_tmp_175;
  wire mux_tmp_393;
  wire mux_tmp_395;
  wire mux_tmp_399;
  wire and_tmp_35;
  wire or_tmp_497;
  wire mux_tmp_405;
  wire not_tmp_236;
  wire mux_tmp_418;
  wire nand_tmp_52;
  wire or_tmp_561;
  wire or_tmp_562;
  wire mux_tmp_448;
  wire or_tmp_566;
  wire mux_tmp_450;
  wire mux_tmp_452;
  wire mux_tmp_456;
  wire mux_tmp_457;
  wire not_tmp_249;
  wire or_tmp_574;
  wire nand_tmp_59;
  wire or_tmp_577;
  wire mux_tmp_458;
  wire mux_tmp_460;
  wire mux_tmp_462;
  wire nand_tmp_62;
  wire mux_tmp_481;
  wire mux_tmp_483;
  wire mux_tmp_484;
  wire mux_tmp_485;
  wire mux_tmp_486;
  wire nand_tmp_65;
  wire nand_tmp_66;
  wire mux_tmp_501;
  wire mux_tmp_502;
  wire or_tmp_604;
  wire mux_tmp_505;
  wire nand_tmp_70;
  wire and_tmp_51;
  wire and_tmp_52;
  wire mux_tmp_518;
  wire mux_tmp_522;
  wire mux_tmp_575;
  wire mux_tmp_581;
  wire not_tmp_280;
  wire or_tmp_695;
  wire mux_tmp_583;
  wire or_tmp_703;
  wire or_tmp_704;
  wire mux_tmp_589;
  wire mux_tmp_591;
  wire mux_tmp_593;
  wire mux_tmp_597;
  wire and_dcpl_821;
  wire and_dcpl_831;
  wire nor_tmp_291;
  wire mux_tmp_604;
  wire or_tmp_723;
  wire or_tmp_724;
  wire mux_tmp_612;
  wire mux_tmp_614;
  wire or_dcpl_209;
  wire or_dcpl_263;
  wire and_tmp_58;
  wire or_tmp_853;
  wire and_tmp_61;
  wire and_tmp_64;
  wire and_tmp_67;
  wire and_tmp_70;
  wire and_tmp_73;
  wire and_tmp_75;
  wire and_tmp_77;
  wire and_tmp_80;
  wire and_tmp_83;
  wire and_tmp_86;
  wire and_tmp_89;
  wire and_tmp_92;
  wire and_tmp_95;
  wire and_tmp_98;
  wire and_tmp_101;
  wire and_tmp_104;
  wire and_tmp_107;
  wire and_tmp_110;
  wire and_tmp_113;
  wire and_tmp_116;
  wire and_tmp_119;
  wire and_tmp_121;
  wire and_tmp_123;
  wire and_tmp_126;
  wire and_tmp_129;
  wire and_tmp_132;
  wire and_tmp_135;
  wire and_tmp_138;
  wire and_tmp_141;
  wire and_tmp_144;
  wire and_tmp_147;
  wire and_tmp_150;
  wire and_tmp_153;
  wire and_tmp_156;
  wire and_tmp_159;
  wire and_tmp_162;
  wire and_tmp_165;
  wire and_tmp_167;
  wire and_tmp_169;
  wire and_tmp_172;
  wire and_tmp_175;
  wire and_tmp_178;
  wire and_tmp_181;
  wire and_tmp_184;
  wire and_tmp_187;
  wire and_tmp_190;
  wire and_tmp_193;
  wire and_tmp_196;
  wire and_tmp_199;
  wire and_tmp_202;
  wire and_tmp_205;
  wire and_tmp_208;
  wire and_tmp_211;
  wire and_tmp_213;
  wire and_tmp_215;
  wire and_tmp_218;
  wire and_tmp_221;
  wire and_tmp_224;
  wire and_tmp_227;
  wire and_tmp_230;
  wire and_tmp_233;
  wire and_tmp_236;
  wire and_tmp_239;
  wire and_tmp_242;
  wire and_tmp_245;
  wire and_tmp_248;
  wire and_tmp_251;
  wire and_tmp_254;
  wire and_tmp_257;
  wire and_tmp_259;
  wire and_tmp_261;
  wire and_tmp_264;
  wire and_tmp_267;
  wire and_tmp_270;
  wire and_tmp_273;
  wire and_tmp_276;
  wire and_tmp_279;
  wire and_tmp_282;
  wire and_tmp_285;
  wire and_tmp_288;
  wire and_tmp_291;
  wire and_tmp_294;
  wire and_tmp_297;
  wire and_tmp_300;
  wire and_tmp_303;
  wire and_tmp_305;
  wire and_tmp_307;
  wire and_tmp_310;
  wire and_tmp_313;
  wire and_tmp_316;
  wire and_tmp_319;
  wire and_tmp_322;
  wire and_tmp_325;
  wire and_tmp_328;
  wire and_tmp_331;
  wire and_tmp_334;
  wire and_tmp_337;
  wire and_tmp_340;
  wire and_tmp_343;
  wire and_tmp_346;
  wire and_tmp_349;
  wire and_tmp_351;
  wire and_tmp_353;
  wire and_tmp_356;
  wire and_tmp_359;
  wire and_tmp_362;
  wire and_tmp_365;
  wire and_tmp_368;
  wire and_tmp_371;
  wire and_tmp_374;
  wire and_tmp_377;
  wire and_tmp_380;
  wire and_tmp_383;
  wire and_tmp_386;
  wire and_tmp_389;
  wire and_tmp_392;
  wire and_tmp_395;
  wire and_tmp_397;
  wire and_tmp_399;
  wire and_tmp_402;
  wire and_tmp_405;
  wire and_tmp_408;
  wire and_tmp_411;
  wire and_tmp_414;
  wire and_tmp_417;
  wire or_tmp_1480;
  wire or_tmp_1481;
  wire or_tmp_2017;
  wire or_tmp_2027;
  wire or_tmp_2033;
  wire or_tmp_2041;
  wire or_tmp_2056;
  wire or_tmp_2094;
  wire or_tmp_2314;
  wire or_tmp_2315;
  wire or_tmp_2337;
  wire or_tmp_2350;
  wire or_tmp_2354;
  wire exit_LOAD_LOOP_lpi_2_dfm_4;
  wire exit_LOAD_LOOP_for_lpi_2_dfm_3_mx0w0;
  wire exit_LOAD_LOOP_sva_3;
  wire exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_3;
  wire LOAD_LOOP_for_if_2_for_equal_tmp_2_mx0w0;
  wire exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_mx0w0;
  wire exit_LOAD_LOOP_for_if_for_sva_1_mx0w0;
  wire [2:0] LOAD_LOOP_for_if_for_m_2_0_lpi_2_mx1;
  wire LOAD_LOOP_for_if_for_for_if_nor_cse_sva_1;
  wire exit_LOAD_LOOP_for_if_for_for_sva_mx0w0;
  wire exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0;
  wire [2:0] LOAD_LOOP_for_print_buf_lpi_2_mx2_7_5;
  wire lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1;
  reg lfst_exit_LOAD_LOOP_for_1_lpi_2;
  reg lfst_exit_LOAD_LOOP_sva;
  wire lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2_mx0w0;
  wire [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0_mx0w0;
  reg lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2;
  reg lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2;
  reg LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
  reg LOAD_LOOP_for_if_2_for_or_tmp_1;
  wire LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  wire LOAD_LOOP_for_if_2_for_and_181_cse_1;
  reg exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_1;
  reg LOAD_LOOP_for_if_2_for_equal_tmp_1;
  reg LOAD_LOOP_for_if_2_for_mux_11_itm_1;
  reg LOAD_LOOP_for_if_2_for_equal_tmp_1_1;
  reg exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_1;
  reg exit_LOAD_LOOP_for_if_2_for_sva_1_1;
  reg exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_1;
  reg exit_LOAD_LOOP_for_if_for_sva_1_1;
  reg [7:0] LOAD_LOOP_for_print_buf_lpi_2;
  reg [7:0] LOAD_LOOP_for_print_buf_sva_1_1;
  wire [8:0] nl_LOAD_LOOP_for_print_buf_sva_1_1;
  reg LOAD_LOOP_for_if_2_for_nor_tmp_1;
  wire LOAD_LOOP_for_if_2_for_and_180_cse_1;
  wire LOAD_LOOP_for_if_2_for_for_and_250_tmp_1;
  wire exitL_exit_LOAD_CTRL_LOOP2_lpi_2_dfm_1;
  reg LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_16_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_0_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_15_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_1_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_14_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_2_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_13_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_3_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_12_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_4_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_11_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_5_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_10_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_6_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_9_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_7_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_4_8_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_15_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_1_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_14_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_2_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_13_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_3_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_12_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_4_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_11_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_5_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_10_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_6_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_9_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_7_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_8_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_3_0_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_1_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_2_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_3_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_4_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_5_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_6_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_7_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_2_0_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_1_1_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_1_2_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_1_3_sva_1;
  wire LOAD_LOOP_for_if_for_for_and_stg_1_0_sva_1;
  reg LOAD_LOOP_for_asn_6_itm_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_61_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_0_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_60_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_1_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_59_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_2_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_58_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_3_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_57_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_4_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_56_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_5_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_55_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_6_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_54_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_7_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_53_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_8_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_52_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_9_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_51_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_10_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_50_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_11_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_49_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_12_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_48_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_13_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_47_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_14_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_46_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_15_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_45_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_16_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_44_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_17_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_43_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_18_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_42_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_19_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_41_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_20_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_40_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_21_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_39_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_22_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_38_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_23_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_37_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_24_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_36_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_25_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_35_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_26_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_34_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_27_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_33_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_28_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_32_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_29_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_31_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_5_30_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_31_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_30_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_0_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_1_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_2_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_3_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_4_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_5_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_6_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_7_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_8_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_9_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_10_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_11_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_12_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_13_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_14_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_15_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_16_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_17_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_18_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_19_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_20_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_21_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_22_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_23_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_24_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_25_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_26_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_27_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_28_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_4_29_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_14_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_15_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_0_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_1_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_2_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_3_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_4_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_5_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_6_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_7_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_8_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_9_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_10_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_11_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_12_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_3_13_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_6_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_7_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_0_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_1_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_2_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_3_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_4_sva_1;
  wire LOAD_LOOP_for_if_2_for_for_and_stg_2_5_sva_1;
  reg LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1;
  reg LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1;
  reg LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1;
  reg LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1;
  reg LOAD_LOOP_for_if_2_for_for_asn_itm_2;
  reg lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2;
  reg LOAD_BATCH_LOOP_stage_v_2;
  reg exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2;
  reg LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3;
  reg exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3;
  reg lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2;
  reg [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0;
  reg LOAD_BATCH_LOOP_stage_v_3;
  reg [4:0] LOAD_LOOP_fl_5_0_sva_4_0;
  reg [231:0] conf_info_crt_sva_231_0;
  wire [2:0] LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_mx1;
  wire LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_and_cse_1;
  wire LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_nor_1_cse_1;
  wire LOAD_LOOP_for_if_2_for_equal_tmp_mx0w0;
  wire LOAD_LOOP_for_if_2_for_equal_tmp_1_mx0w0;
  wire lfst_exit_LOAD_LOOP_sva_dfm_1_mx0w1;
  wire [3:0] LOAD_LOOP_for_if_2_for_for_acc_2_psp_1;
  wire [4:0] nl_LOAD_LOOP_for_if_2_for_for_acc_2_psp_1;
  wire [2:0] LOAD_LOOP_for_if_2_for_for_row_norm_2_0_lpi_2_dfm_1;
  reg [4:0] LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2;
  reg [4:0] LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_1;
  reg [4:0] LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_2_1;
  reg exit_LOAD_LOOP_for_if_2_for_for_sva_1;
  wire LOAD_LOOP_for_if_2_for_and_178_m1c_1;
  reg exit_LOAD_LOOP_for_lpi_2_dfm_3;
  reg lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2;
  reg [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0;
  reg LOAD_LOOP_for_asn_2_itm_1;
  reg exit_LOAD_LOOP_for_if_for_for_sva_1;
  reg LOAD_LOOP_for_if_2_for_for_asn_itm_1;
  reg LOAD_BATCH_LOOP_stage_0_3;
  reg [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0;
  reg LOAD_BATCH_LOOP_stage_0_2;
  reg [2:0] LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_5_3;
  reg [2:0] LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0;
  reg LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1;
  reg exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_1;
  reg LOAD_BATCH_LOOP_asn_itm_1;
  reg LOAD_LOOP_for_if_2_for_for_asn_126_itm_2;
  reg LOAD_BATCH_LOOP_asn_itm_2;
  reg LOAD_LOOP_for_if_2_for_equal_tmp_2_2;
  reg [2:0] LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3;
  reg [1:0] LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1;
  reg exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_2;
  reg LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_2;
  reg LOAD_BATCH_LOOP_stage_0_1;
  reg LOAD_BATCH_LOOP_stage_0;
  reg [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0;
  reg lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2;
  reg exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  reg exitL_exit_LOAD_LOOP_for_if_2_for_sva_1;
  reg LOAD_LOOP_for_asn_sft_lpi_2;
  reg sfi_operator_8_false_operator_8_false_nor_cse_lpi_2;
  reg [5:0] LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1;
  wire [6:0] nl_LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1;
  reg exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_1;
  reg operator_8_false_operator_8_false_nor_cse_lpi_2;
  reg LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st_1;
  reg LOAD_BATCH_LOOP_stage_v;
  reg LOAD_LOOP_for_if_for_for_and_108_psp;
  reg LOAD_LOOP_for_if_for_for_and_107_psp;
  reg LOAD_LOOP_for_if_for_for_and_106_psp;
  reg LOAD_LOOP_for_if_for_for_and_105_psp;
  reg LOAD_LOOP_for_if_for_for_and_104_psp;
  reg LOAD_LOOP_for_if_for_for_and_103_psp;
  reg LOAD_LOOP_for_if_for_for_and_102_psp;
  reg LOAD_LOOP_for_if_for_for_and_101_psp;
  reg LOAD_LOOP_for_if_for_for_and_100_psp;
  reg LOAD_LOOP_for_if_for_for_and_99_psp;
  reg LOAD_LOOP_for_if_for_for_and_98_psp;
  reg LOAD_LOOP_for_if_for_for_and_97_psp;
  reg LOAD_LOOP_for_if_for_for_and_96_psp;
  reg LOAD_LOOP_for_if_for_for_and_95_psp;
  reg LOAD_LOOP_for_if_for_for_and_94_psp;
  reg LOAD_LOOP_for_if_for_for_and_93_psp;
  reg LOAD_LOOP_for_if_for_for_and_92_psp;
  reg LOAD_LOOP_for_if_for_for_and_91_psp;
  reg LOAD_LOOP_for_if_for_for_and_90_psp;
  reg LOAD_LOOP_for_if_for_for_and_89_psp;
  reg LOAD_LOOP_for_if_for_for_and_88_psp;
  reg LOAD_LOOP_for_if_for_for_and_87_psp;
  reg LOAD_LOOP_for_if_for_for_and_86_psp;
  reg LOAD_LOOP_for_if_for_for_and_85_psp;
  reg LOAD_LOOP_for_if_for_for_and_84_psp;
  reg LOAD_LOOP_for_if_for_for_and_83_psp;
  reg LOAD_LOOP_for_if_for_for_and_82_psp;
  reg LOAD_LOOP_for_if_for_for_and_81_psp;
  reg LOAD_LOOP_for_if_for_for_and_80_psp;
  reg LOAD_LOOP_for_if_for_for_and_79_psp;
  reg LOAD_LOOP_for_if_for_for_and_78_psp;
  reg LOAD_LOOP_for_if_for_for_and_77_psp;
  reg LOAD_LOOP_for_if_for_for_and_76_psp;
  reg LOAD_LOOP_for_if_for_for_and_75_psp;
  reg LOAD_LOOP_for_if_for_for_and_74_psp;
  reg LOAD_LOOP_for_if_for_for_and_73_psp;
  reg LOAD_LOOP_for_if_for_for_and_72_psp;
  reg LOAD_LOOP_for_if_for_for_and_71_psp;
  reg LOAD_LOOP_for_if_for_for_and_70_psp;
  reg LOAD_LOOP_for_if_for_for_and_69_psp;
  reg LOAD_LOOP_for_if_for_for_and_68_psp;
  reg LOAD_LOOP_for_if_for_for_and_67_psp;
  reg LOAD_LOOP_for_if_for_for_and_66_psp;
  reg LOAD_LOOP_for_if_for_for_and_65_psp;
  reg LOAD_LOOP_for_if_for_for_and_64_psp;
  reg LOAD_LOOP_for_if_for_for_and_63_psp;
  reg LOAD_LOOP_for_if_for_for_and_62_psp;
  reg LOAD_LOOP_for_if_for_for_and_61_psp;
  reg LOAD_LOOP_for_if_for_for_and_60_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_249_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_248_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_247_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_246_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_245_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_244_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_243_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_242_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_241_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_240_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_239_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_238_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_237_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_236_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_235_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_234_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_233_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_232_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_231_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_230_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_229_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_228_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_227_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_226_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_225_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_224_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_223_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_222_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_221_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_220_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_219_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_218_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_217_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_216_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_215_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_214_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_213_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_212_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_211_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_210_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_209_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_208_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_207_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_206_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_205_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_204_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_203_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_202_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_201_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_200_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_199_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_198_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_197_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_196_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_195_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_194_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_193_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_192_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_191_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_190_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_189_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_188_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_187_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_186_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_185_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_184_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_183_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_182_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_181_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_180_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_179_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_178_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_177_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_176_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_175_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_174_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_173_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_172_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_171_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_170_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_169_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_168_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_167_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_166_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_165_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_164_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_163_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_162_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_161_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_160_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_159_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_158_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_157_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_156_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_155_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_154_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_153_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_152_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_151_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_150_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_149_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_148_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_147_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_146_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_145_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_144_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_143_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_142_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_141_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_140_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_139_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_138_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_137_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_136_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_135_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_134_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_133_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_132_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_131_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_130_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_129_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_128_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_127_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_126_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_125_psp;
  reg LOAD_LOOP_for_if_2_for_for_and_124_psp;
  wire [2:0] LOAD_LOOP_for_if_for_m_2_0_sva_1_mx0w1;
  wire [3:0] nl_LOAD_LOOP_for_if_for_m_2_0_sva_1_mx0w1;
  wire exit_LOAD_LOOP_lpi_2_dfm_1_mx0w0;
  reg exit_LOAD_LOOP_lpi_2_dfm_1;
  wire exit_LOAD_LOOP_for_if_for_lpi_2_dfm_mx0w0;
  reg exit_LOAD_LOOP_for_if_for_lpi_2_dfm;
  reg exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm;
  wire [4:0] LOAD_LOOP_for_print_buf_lpi_2_mx1_4_0;
  wire exitL_exit_LOAD_LOOP_for_if_2_for_sva_1_mx0w0;
  wire [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1;
  wire exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1;
  wire or_1873_tmp;
  wire and_1304_tmp;
  reg reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse;
  reg reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse;
  reg reg_done_rsci_ivld_core_psct_cse;
  reg reg_dma_read_chnl_rsci_irdy_core_psct_cse;
  reg reg_dma_read_ctrl_rsci_ivld_core_psct_cse;
  reg reg_plm_kernel_rsci_ivld_core_psct_cse;
  reg reg_buf_linear_rsci_ivld_core_psct_cse;
  reg reg_conf_info_rsci_irdy_core_psct_cse;
  wire LOAD_LOOP_for_if_for_and_cse;
  wire LOAD_LOOP_for_if_2_for_if_and_128_cse;
  wire LOAD_LOOP_for_if_for_and_2_cse;
  wire LOAD_LOOP_for_if_for_and_3_cse;
  wire LOAD_LOOP_for_if_for_for_and_111_cse;
  wire and_3195_cse;
  wire nor_752_cse;
  wire LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse;
  wire LOAD_LOOP_for_and_2_cse;
  wire LOAD_LOOP_for_if_2_for_for_and_259_cse;
  wire LOAD_LOOP_for_if_2_for_and_205_cse;
  wire LOAD_LOOP_for_if_2_for_for_and_257_cse;
  wire operator_8_false_and_cse;
  wire or_654_cse;
  wire LOAD_LOOP_for_if_for_for_n_and_1_cse;
  wire LOAD_LOOP_fl_and_cse;
  wire LOAD_LOOP_for_and_5_cse;
  wire or_941_cse;
  wire or_939_cse;
  wire or_967_cse;
  wire nor_307_cse;
  wire or_960_cse;
  wire nor_304_cse;
  wire nor_302_cse;
  wire or_950_cse;
  wire and_3220_cse;
  wire nand_222_cse;
  wire nand_213_cse;
  wire nand_195_cse;
  wire or_810_cse;
  wire and_3197_cse;
  wire or_9_cse;
  wire or_75_cse;
  wire nor_32_cse;
  wire or_44_cse;
  wire and_3266_cse;
  wire or_750_cse;
  wire or_755_cse;
  wire LOAD_LOOP_for_LOAD_LOOP_nand_cse;
  wire nor_37_cse;
  wire or_93_cse;
  wire and_3192_cse;
  wire nor_225_cse;
  wire or_41_cse;
  wire and_3198_cse;
  wire or_42_cse;
  wire nor_566_cse;
  wire or_539_cse;
  wire nor_55_cse;
  wire or_481_cse;
  wire nor_113_cse;
  wire or_631_cse;
  wire or_439_cse;
  wire nor_778_cse;
  wire or_289_cse;
  wire or_305_cse;
  wire or_309_cse;
  wire or_313_cse;
  wire or_317_cse;
  wire or_321_cse;
  wire or_325_cse;
  wire or_329_cse;
  wire or_333_cse;
  wire or_337_cse;
  wire or_341_cse;
  wire or_345_cse;
  wire or_349_cse;
  wire or_353_cse;
  wire or_357_cse;
  wire nand_106_cse;
  wire or_365_cse;
  wire or_373_cse;
  wire or_377_cse;
  wire or_381_cse;
  wire or_385_cse;
  wire or_389_cse;
  wire or_393_cse;
  wire nand_102_cse;
  wire or_401_cse;
  wire or_409_cse;
  wire or_413_cse;
  wire or_417_cse;
  wire or_421_cse;
  wire or_429_cse;
  wire or_632_cse;
  wire [4:0] LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1;
  wire or_2860_cse;
  wire or_513_cse;
  wire nand_223_cse;
  wire nand_224_cse;
  wire nand_225_cse;
  wire nand_212_cse;
  wire nand_214_cse;
  wire nand_215_cse;
  wire nand_218_cse;
  wire nand_194_cse;
  wire nand_196_cse;
  wire nand_197_cse;
  wire nand_199_cse;
  wire nand_163_cse;
  wire nand_164_cse;
  wire nand_165_cse;
  wire nand_167_cse;
  wire or_101_cse;
  wire mux_335_cse;
  wire mux_107_cse;
  wire or_634_cse;
  wire mux_491_cse;
  wire mux_497_cse;
  wire mux_510_cse;
  wire or_843_cse;
  wire mux_609_cse;
  wire mux_619_cse;
  wire mux_575_cse;
  wire or_588_cse;
  wire or_771_cse;
  wire LOAD_LOOP_for_and_9_cse;
  wire and_834_cse;
  wire nand_24_cse;
  wire or_197_cse;
  wire mux_481_cse;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d_reg;
  wire [31:0] LOAD_LOOP_for_if_2_for_for_if_mux_rmff;
  reg [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d_reg;
  wire [13:0] LOAD_LOOP_for_if_2_for_for_else_index_in_mux_rmff;
  reg [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d_reg;
  wire [13:0] LOAD_LOOP_for_if_2_for_for_if_index_in_mux_rmff;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_iff;
  wire and_2372_rmff;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_2370_rmff;
  wire or_dcpl_395;
  wire or_dcpl_401;
  wire LOAD_LOOP_for_if_for_for_and_tmp_1;
  wire LOAD_LOOP_for_if_2_for_for_and_251_tmp_1;
  wire or_2901_tmp;
  wire or_2899_tmp;
  wire LOAD_LOOP_for_if_2_for_and_191_tmp;
  wire or_2895_tmp;
  wire or_2893_tmp;
  wire LOAD_LOOP_for_if_2_for_and_187_tmp;
  wire LOAD_LOOP_for_if_2_for_and_176_m1c_1;
  wire LOAD_LOOP_for_if_2_for_and_199_cse;
  wire or_461_itm;
  wire mux_612_itm;
  wire [13:0] z_out_1;
  wire [20:0] nl_z_out_1;
  wire mux_tmp;
  wire [16:0] z_out_4;
  wire signed [22:0] nl_z_out_4;
  wire [15:0] z_out_5;
  wire [23:0] nl_z_out_5;
  wire [15:0] z_out_6;
  wire [23:0] nl_z_out_6;
  wire [2:0] z_out_7;
  wire [2:0] z_out_8;
  wire or_tmp_2431;
  wire [2:0] z_out_9;
  wire [3:0] nl_z_out_9;
  wire [16:0] z_out_10;
  wire [17:0] nl_z_out_10;
  wire [8:0] z_out_11;
  wire [15:0] z_out_12;
  wire [16:0] nl_z_out_12;
  wire [8:0] z_out_13;
  wire [9:0] nl_z_out_13;
  reg [15:0] LOAD_LOOP_for_mul_cse_lpi_2;
  reg [15:0] LOAD_LOOP_for_ac_int_cctor_lpi_2;
  reg [2:0] LOAD_LOOP_for_if_for_m_2_0_lpi_2;
  reg [2:0] LOAD_LOOP_for_if_for_for_n_2_0_lpi_2;
  reg [15:0] LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2;
  reg [4:0] LOAD_LOOP_for_if_2_for_row_4_0_lpi_2;
  reg [7:0] pad_sva;
  reg [6:0] n_w_in_acc_psp_sva;
  wire [7:0] nl_n_w_in_acc_psp_sva;
  reg [6:0] n_h_in_acc_psp_sva;
  wire [7:0] nl_n_h_in_acc_psp_sva;
  reg [15:0] batch_size_mul_4_cse_sva;
  reg [15:0] batch_size_mul_3_cse_sva;
  reg [15:0] batch_size_mul_2_cse_sva;
  reg [15:0] batch_size_mul_1_cse_sva;
  reg [15:0] batch_size_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_24_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_23_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_25_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_22_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_26_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_21_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_27_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_20_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_28_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_19_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_29_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_18_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_30_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_17_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_31_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_32_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_33_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_34_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_35_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_36_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_37_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_38_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_39_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_40_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_41_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_42_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_43_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_44_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_45_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_46_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_47_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_plm_tmp_f_data_48_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_3_17_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_17_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_2_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_4_17_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_17_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_1_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_5_17_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_17_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_8_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_9_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_7_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_10_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_6_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_11_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_5_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_12_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_4_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_13_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_3_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_14_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_2_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_15_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_1_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_16_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_0_0_sva;
  reg [31:0] LOAD_BATCH_LOOP_buf_tmp_lin_data_6_17_sva;
  reg [7:0] LOAD_LOOP_for_print_buf_lpi_2_dfm_3;
  reg [15:0] LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2;
  reg operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1;
  reg [2:0] LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3;
  reg [2:0] LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4;
  reg [4:0] LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3;
  reg [4:0] LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4;
  reg LOAD_LOOP_for_asn_sft_lpi_2_dfm_1;
  reg sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1;
  reg LOAD_BATCH_LOOP_stage_v_1;
  reg exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st;
  reg LOAD_LOOP_for_asn_2_itm;
  reg LOAD_LOOP_for_if_2_for_for_asn_itm;
  reg LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st;
  reg exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st;
  reg LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st;
  reg [4:0] LOAD_LOOP_for_if_2_for_row_4_0_sva_1_1;
  reg [31:0] LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1;
  reg [2:0] LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_2_1;
  reg [2:0] LOAD_LOOP_for_if_for_m_2_0_sva_1_1;
  reg [2:0] LOAD_LOOP_for_if_for_for_n_2_0_sva_1_1;
  reg LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_1;
  reg [13:0] LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1;
  wire [14:0] nl_LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1;
  reg [4:0] LOAD_LOOP_for_k_5_0_lpi_2_4_0;
  reg [3:0] LOAD_BATCH_LOOP_b_4_0_sva_3_0;
  reg [2:0] LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3;
  reg [2:0] LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_0;
  reg lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2;
  reg [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0;
  reg [1:0] lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_1_0;
  wire dma_read_ctrl_rsci_idat_15_0_mx0c2;
  wire dma_read_ctrl_rsci_idat_47_32_mx0c1;
  wire plm_kernel_rsci_idat_31_0_mx0c1;
  wire plm_kernel_rsci_idat_63_32_mx0c1;
  wire plm_kernel_rsci_idat_95_64_mx0c1;
  wire plm_kernel_rsci_idat_127_96_mx0c1;
  wire plm_kernel_rsci_idat_159_128_mx0c1;
  wire plm_kernel_rsci_idat_191_160_mx0c1;
  wire plm_kernel_rsci_idat_223_192_mx0c1;
  wire plm_kernel_rsci_idat_255_224_mx0c1;
  wire plm_kernel_rsci_idat_287_256_mx0c1;
  wire plm_kernel_rsci_idat_319_288_mx0c1;
  wire plm_kernel_rsci_idat_351_320_mx0c1;
  wire plm_kernel_rsci_idat_383_352_mx0c1;
  wire plm_kernel_rsci_idat_415_384_mx0c1;
  wire plm_kernel_rsci_idat_447_416_mx0c1;
  wire plm_kernel_rsci_idat_479_448_mx0c1;
  wire plm_kernel_rsci_idat_511_480_mx0c1;
  wire plm_kernel_rsci_idat_543_512_mx0c1;
  wire plm_kernel_rsci_idat_575_544_mx0c1;
  wire plm_kernel_rsci_idat_607_576_mx0c1;
  wire plm_kernel_rsci_idat_639_608_mx0c1;
  wire plm_kernel_rsci_idat_671_640_mx0c1;
  wire plm_kernel_rsci_idat_703_672_mx0c1;
  wire plm_kernel_rsci_idat_735_704_mx0c1;
  wire plm_kernel_rsci_idat_767_736_mx0c1;
  wire plm_kernel_rsci_idat_799_768_mx0c1;
  wire plm_kernel_rsci_idat_831_800_mx0c1;
  wire plm_kernel_rsci_idat_863_832_mx0c1;
  wire plm_kernel_rsci_idat_895_864_mx0c1;
  wire plm_kernel_rsci_idat_927_896_mx0c1;
  wire plm_kernel_rsci_idat_959_928_mx0c1;
  wire plm_kernel_rsci_idat_991_960_mx0c1;
  wire plm_kernel_rsci_idat_1023_992_mx0c1;
  wire plm_kernel_rsci_idat_1055_1024_mx0c1;
  wire plm_kernel_rsci_idat_1087_1056_mx0c1;
  wire plm_kernel_rsci_idat_1119_1088_mx0c1;
  wire plm_kernel_rsci_idat_1151_1120_mx0c1;
  wire plm_kernel_rsci_idat_1183_1152_mx0c1;
  wire plm_kernel_rsci_idat_1215_1184_mx0c1;
  wire plm_kernel_rsci_idat_1247_1216_mx0c1;
  wire plm_kernel_rsci_idat_1279_1248_mx0c1;
  wire plm_kernel_rsci_idat_1311_1280_mx0c1;
  wire plm_kernel_rsci_idat_1343_1312_mx0c1;
  wire plm_kernel_rsci_idat_1375_1344_mx0c1;
  wire plm_kernel_rsci_idat_1407_1376_mx0c1;
  wire plm_kernel_rsci_idat_1439_1408_mx0c1;
  wire plm_kernel_rsci_idat_1471_1440_mx0c1;
  wire plm_kernel_rsci_idat_1503_1472_mx0c1;
  wire plm_kernel_rsci_idat_1535_1504_mx0c1;
  wire plm_kernel_rsci_idat_1567_1536_mx0c1;
  wire buf_linear_rsci_idat_31_0_mx0c1;
  wire buf_linear_rsci_idat_63_32_mx0c1;
  wire buf_linear_rsci_idat_95_64_mx0c1;
  wire buf_linear_rsci_idat_127_96_mx0c1;
  wire buf_linear_rsci_idat_159_128_mx0c1;
  wire buf_linear_rsci_idat_191_160_mx0c1;
  wire buf_linear_rsci_idat_223_192_mx0c1;
  wire buf_linear_rsci_idat_255_224_mx0c1;
  wire buf_linear_rsci_idat_287_256_mx0c1;
  wire buf_linear_rsci_idat_319_288_mx0c1;
  wire buf_linear_rsci_idat_351_320_mx0c1;
  wire buf_linear_rsci_idat_383_352_mx0c1;
  wire buf_linear_rsci_idat_415_384_mx0c1;
  wire buf_linear_rsci_idat_447_416_mx0c1;
  wire buf_linear_rsci_idat_479_448_mx0c1;
  wire buf_linear_rsci_idat_511_480_mx0c1;
  wire buf_linear_rsci_idat_543_512_mx0c1;
  wire buf_linear_rsci_idat_575_544_mx0c1;
  wire buf_linear_rsci_idat_607_576_mx0c1;
  wire buf_linear_rsci_idat_639_608_mx0c1;
  wire buf_linear_rsci_idat_671_640_mx0c1;
  wire buf_linear_rsci_idat_703_672_mx0c1;
  wire buf_linear_rsci_idat_735_704_mx0c1;
  wire buf_linear_rsci_idat_767_736_mx0c1;
  wire buf_linear_rsci_idat_799_768_mx0c1;
  wire buf_linear_rsci_idat_831_800_mx0c1;
  wire buf_linear_rsci_idat_863_832_mx0c1;
  wire buf_linear_rsci_idat_895_864_mx0c1;
  wire buf_linear_rsci_idat_927_896_mx0c1;
  wire buf_linear_rsci_idat_959_928_mx0c1;
  wire buf_linear_rsci_idat_991_960_mx0c1;
  wire buf_linear_rsci_idat_1023_992_mx0c1;
  wire buf_linear_rsci_idat_1055_1024_mx0c1;
  wire buf_linear_rsci_idat_1087_1056_mx0c1;
  wire buf_linear_rsci_idat_1119_1088_mx0c1;
  wire buf_linear_rsci_idat_1151_1120_mx0c1;
  wire buf_linear_rsci_idat_1183_1152_mx0c1;
  wire buf_linear_rsci_idat_1215_1184_mx0c1;
  wire buf_linear_rsci_idat_1247_1216_mx0c1;
  wire buf_linear_rsci_idat_1279_1248_mx0c1;
  wire buf_linear_rsci_idat_1311_1280_mx0c1;
  wire buf_linear_rsci_idat_1343_1312_mx0c1;
  wire buf_linear_rsci_idat_1375_1344_mx0c1;
  wire buf_linear_rsci_idat_1407_1376_mx0c1;
  wire buf_linear_rsci_idat_1439_1408_mx0c1;
  wire buf_linear_rsci_idat_1471_1440_mx0c1;
  wire buf_linear_rsci_idat_1503_1472_mx0c1;
  wire buf_linear_rsci_idat_1535_1504_mx0c1;
  wire buf_linear_rsci_idat_1567_1536_mx0c1;
  wire buf_linear_rsci_idat_1599_1568_mx0c1;
  wire buf_linear_rsci_idat_1631_1600_mx0c1;
  wire buf_linear_rsci_idat_1663_1632_mx0c1;
  wire buf_linear_rsci_idat_1695_1664_mx0c1;
  wire buf_linear_rsci_idat_1727_1696_mx0c1;
  wire buf_linear_rsci_idat_1759_1728_mx0c1;
  wire buf_linear_rsci_idat_1791_1760_mx0c1;
  wire buf_linear_rsci_idat_1823_1792_mx0c1;
  wire buf_linear_rsci_idat_1855_1824_mx0c1;
  wire buf_linear_rsci_idat_1887_1856_mx0c1;
  wire buf_linear_rsci_idat_1919_1888_mx0c1;
  wire buf_linear_rsci_idat_1951_1920_mx0c1;
  wire buf_linear_rsci_idat_1983_1952_mx0c1;
  wire buf_linear_rsci_idat_2015_1984_mx0c1;
  wire buf_linear_rsci_idat_2047_2016_mx0c1;
  wire buf_linear_rsci_idat_2079_2048_mx0c1;
  wire buf_linear_rsci_idat_2111_2080_mx0c1;
  wire buf_linear_rsci_idat_2143_2112_mx0c1;
  wire buf_linear_rsci_idat_2175_2144_mx0c1;
  wire buf_linear_rsci_idat_2207_2176_mx0c1;
  wire buf_linear_rsci_idat_2239_2208_mx0c1;
  wire buf_linear_rsci_idat_2271_2240_mx0c1;
  wire buf_linear_rsci_idat_2303_2272_mx0c1;
  wire buf_linear_rsci_idat_2335_2304_mx0c1;
  wire buf_linear_rsci_idat_2367_2336_mx0c1;
  wire buf_linear_rsci_idat_2399_2368_mx0c1;
  wire buf_linear_rsci_idat_2431_2400_mx0c1;
  wire buf_linear_rsci_idat_2463_2432_mx0c1;
  wire buf_linear_rsci_idat_2495_2464_mx0c1;
  wire buf_linear_rsci_idat_2527_2496_mx0c1;
  wire buf_linear_rsci_idat_2559_2528_mx0c1;
  wire buf_linear_rsci_idat_2591_2560_mx0c1;
  wire buf_linear_rsci_idat_2623_2592_mx0c1;
  wire buf_linear_rsci_idat_2655_2624_mx0c1;
  wire buf_linear_rsci_idat_2687_2656_mx0c1;
  wire buf_linear_rsci_idat_2719_2688_mx0c1;
  wire buf_linear_rsci_idat_2751_2720_mx0c1;
  wire buf_linear_rsci_idat_2783_2752_mx0c1;
  wire buf_linear_rsci_idat_2815_2784_mx0c1;
  wire buf_linear_rsci_idat_2847_2816_mx0c1;
  wire buf_linear_rsci_idat_2879_2848_mx0c1;
  wire buf_linear_rsci_idat_2911_2880_mx0c1;
  wire buf_linear_rsci_idat_2943_2912_mx0c1;
  wire buf_linear_rsci_idat_2975_2944_mx0c1;
  wire buf_linear_rsci_idat_3007_2976_mx0c1;
  wire buf_linear_rsci_idat_3039_3008_mx0c1;
  wire buf_linear_rsci_idat_3071_3040_mx0c1;
  wire buf_linear_rsci_idat_3103_3072_mx0c1;
  wire buf_linear_rsci_idat_3135_3104_mx0c1;
  wire buf_linear_rsci_idat_3167_3136_mx0c1;
  wire buf_linear_rsci_idat_3199_3168_mx0c1;
  wire buf_linear_rsci_idat_3231_3200_mx0c1;
  wire buf_linear_rsci_idat_3263_3232_mx0c1;
  wire buf_linear_rsci_idat_3295_3264_mx0c1;
  wire buf_linear_rsci_idat_3327_3296_mx0c1;
  wire buf_linear_rsci_idat_3359_3328_mx0c1;
  wire buf_linear_rsci_idat_3391_3360_mx0c1;
  wire buf_linear_rsci_idat_3423_3392_mx0c1;
  wire buf_linear_rsci_idat_3455_3424_mx0c1;
  wire buf_linear_rsci_idat_3487_3456_mx0c1;
  wire buf_linear_rsci_idat_3519_3488_mx0c1;
  wire buf_linear_rsci_idat_3551_3520_mx0c1;
  wire buf_linear_rsci_idat_3583_3552_mx0c1;
  wire buf_linear_rsci_idat_3615_3584_mx0c1;
  wire buf_linear_rsci_idat_3647_3616_mx0c1;
  wire buf_linear_rsci_idat_3679_3648_mx0c1;
  wire buf_linear_rsci_idat_3711_3680_mx0c1;
  wire buf_linear_rsci_idat_3743_3712_mx0c1;
  wire buf_linear_rsci_idat_3775_3744_mx0c1;
  wire buf_linear_rsci_idat_3807_3776_mx0c1;
  wire buf_linear_rsci_idat_3839_3808_mx0c1;
  wire buf_linear_rsci_idat_3871_3840_mx0c1;
  wire buf_linear_rsci_idat_3903_3872_mx0c1;
  wire buf_linear_rsci_idat_3935_3904_mx0c1;
  wire buf_linear_rsci_idat_3967_3936_mx0c1;
  wire buf_linear_rsci_idat_3999_3968_mx0c1;
  wire buf_linear_rsci_idat_4031_4000_mx0c1;
  wire exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0;
  wire [4:0] LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1;
  wire [5:0] nl_LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1;
  wire [4:0] LOAD_LOOP_for_if_2_for_row_4_0_sva_1_mx0w1;
  wire [5:0] nl_LOAD_LOOP_for_if_2_for_row_4_0_sva_1_mx0w1;
  wire [2:0] LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1;
  wire [3:0] nl_LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1;
  wire LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_mx0w0;
  wire LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_mx0w1;
  wire LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1_mx0c1;
  wire [2:0] LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3_mx0w0;
  wire [3:0] nl_LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3_mx0w0;
  wire [2:0] LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3_mx0w0;
  wire [2:0] LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4_mx0w0;
  wire sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1_mx0w0;
  wire LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2_mx0c1;
  wire [7:0] LOAD_LOOP_for_print_buf_lpi_2_dfm_3_mx0w0;
  wire [4:0] LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3_mx0w0;
  wire [4:0] LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4_mx0w0;
  wire LOAD_BATCH_LOOP_stage_v_mx0c0;
  wire LOAD_BATCH_LOOP_stage_v_mx0c1;
  wire LOAD_BATCH_LOOP_stage_v_2_mx0c0;
  wire LOAD_BATCH_LOOP_stage_v_3_mx0c0;
  wire [4:0] LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1;
  wire sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_mx1;
  wire LOAD_LOOP_for_k_5_0_lpi_2_4_0_mx0c1;
  wire LOAD_BATCH_LOOP_stage_v_1_mx0c0;
  wire [31:0] LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_mx0w0;
  wire [31:0] LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
  wire [4:0] LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1;
  wire [8:0] operator_8_false_8_acc_psp_sva_1;
  wire [9:0] nl_operator_8_false_8_acc_psp_sva_1;
  wire [8:0] operator_8_false_5_acc_psp_sva_1;
  wire [9:0] nl_operator_8_false_5_acc_psp_sva_1;
  wire [8:0] operator_8_false_4_acc_psp_sva_1;
  wire [9:0] nl_operator_8_false_4_acc_psp_sva_1;
  wire LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1;
  wire operator_8_false_operator_8_false_nor_cse_sva_1;
  wire [2:0] operator_8_false_1_acc_psp_sva_1;
  wire [4:0] nl_operator_8_false_1_acc_psp_sva_1;
  wire [3:0] operator_8_false_3_acc_psp_sva_1;
  wire [4:0] nl_operator_8_false_3_acc_psp_sva_1;
  wire and_3158_cse;
  wire nor_178_cse;
  wire and_3338_cse;
  wire LOAD_LOOP_for_if_2_for_for_col_and_2_cse;
  wire LOAD_LOOP_for_if_2_for_if_and_132_cse;
  wire and_cse;
  wire and_3316_cse;
  wire and_3318_cse;
  wire mux_1159_itm;
  wire mux_1157_itm;
  wire mux_1158_itm;
  wire operator_8_false_4_acc_itm_3_1;
  wire LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_itm_9_1;
  wire LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_itm_9_1;
  wire operator_8_false_5_acc_itm_4_1;
  wire LOAD_LOOP_for_if_2_for_for_if_aelse_acc_itm_8;
  wire operator_8_false_6_acc_itm_4_1;
  wire [15:0] z_out_15_0;
  wire [15:0] z_out_2_15_0;
  wire [23:0] nl_z_out_2_15_0;
  wire [15:0] z_out_3_15_0;

  wire[0:0] mux_1098_nl;
  wire[0:0] or_1869_nl;
  wire[0:0] LOAD_CTRL_LOOP1_or_nl;
  wire[0:0] LOAD_CTRL_LOOP1_and_2_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] and_808_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] or_2861_nl;
  wire[0:0] or_2862_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] or_452_nl;
  wire[0:0] or_451_nl;
  wire[0:0] or_2868_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] or_474_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] or_467_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] nor_725_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] or_458_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] or_485_nl;
  wire[0:0] or_483_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] or_2436_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] or_538_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] mux_393_nl;
  wire[0:0] and_847_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] and_3196_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] and_849_nl;
  wire[0:0] LOAD_LOOP_for_if_for_LOAD_LOOP_for_if_for_or_1_nl;
  wire[4:0] LOAD_LOOP_for_if_2_for_for_if_1_mux_nl;
  wire[2:0] LOAD_LOOP_for_if_for_for_if_mux_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] nand_48_nl;
  wire[0:0] and_2516_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] and_872_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] and_3194_nl;
  wire[0:0] or_690_nl;
  wire[0:0] mux_420_nl;
  wire[12:0] LOAD_LOOP_for_if_2_for_for_if_index_in_acc_3_nl;
  wire[13:0] nl_LOAD_LOOP_for_if_2_for_for_if_index_in_acc_3_nl;
  wire[12:0] LOAD_LOOP_for_if_2_for_for_if_index_in_mul_7_nl;
  wire[0:0] and_2526_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] and_885_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] mux_473_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] or_749_nl;
  wire[0:0] or_766_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] nand_64_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] and_2666_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] and_899_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] LOAD_LOOP_for_if_for_mux_11_nl;
  wire[0:0] LOAD_LOOP_for_if_for_mux_12_nl;
  wire[4:0] LOAD_LOOP_for_mux_7_nl;
  wire[0:0] LOAD_LOOP_for_and_1_nl;
  wire[0:0] LOAD_BATCH_LOOP_b_not_1_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] LOAD_LOOP_for_k_and_nl;
  wire[0:0] LOAD_LOOP_for_k_and_1_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] nand_269_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] nand_337_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] nand_336_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] nand_268_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] nand_267_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] nand_266_nl;
  wire[0:0] mux_632_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] nand_265_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] nand_264_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] nand_263_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] nand_262_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] nand_261_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] nand_260_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] nand_259_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] nand_258_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] nand_257_nl;
  wire[0:0] mux_653_nl;
  wire[0:0] nand_256_nl;
  wire[0:0] mux_652_nl;
  wire[0:0] mux_655_nl;
  wire[0:0] mux_654_nl;
  wire[0:0] nand_255_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] nand_335_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] nand_334_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] nand_254_nl;
  wire[0:0] mux_663_nl;
  wire[0:0] nand_253_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] nand_252_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] nand_251_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] nand_250_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] nand_249_nl;
  wire[0:0] mux_673_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] nand_248_nl;
  wire[0:0] mux_675_nl;
  wire[0:0] nand_247_nl;
  wire[0:0] mux_674_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] mux_676_nl;
  wire[0:0] nand_246_nl;
  wire[0:0] mux_679_nl;
  wire[0:0] nand_245_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] mux_681_nl;
  wire[0:0] nand_244_nl;
  wire[0:0] mux_680_nl;
  wire[0:0] mux_683_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] nand_243_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] nand_242_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] mux_687_nl;
  wire[0:0] mux_686_nl;
  wire[0:0] nand_241_nl;
  wire[0:0] mux_689_nl;
  wire[0:0] mux_688_nl;
  wire[0:0] nand_333_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] nand_332_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] mux_693_nl;
  wire[0:0] mux_692_nl;
  wire[0:0] nand_240_nl;
  wire[0:0] mux_695_nl;
  wire[0:0] nand_239_nl;
  wire[0:0] mux_694_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] nand_238_nl;
  wire[0:0] mux_696_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] nand_237_nl;
  wire[0:0] mux_701_nl;
  wire[0:0] nand_236_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] mux_703_nl;
  wire[0:0] mux_702_nl;
  wire[0:0] nand_235_nl;
  wire[0:0] mux_705_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] nand_234_nl;
  wire[0:0] mux_707_nl;
  wire[0:0] nand_233_nl;
  wire[0:0] mux_706_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] nand_232_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] nand_231_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] mux_713_nl;
  wire[0:0] nand_230_nl;
  wire[0:0] mux_712_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] mux_714_nl;
  wire[0:0] nand_229_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] nand_228_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] mux_718_nl;
  wire[0:0] nand_227_nl;
  wire[0:0] mux_722_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] mux_720_nl;
  wire[0:0] and_944_nl;
  wire[0:0] and_943_nl;
  wire[0:0] mux_725_nl;
  wire[0:0] mux_724_nl;
  wire[0:0] mux_723_nl;
  wire[0:0] nor_694_nl;
  wire[0:0] and_946_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] mux_727_nl;
  wire[0:0] mux_726_nl;
  wire[0:0] and_950_nl;
  wire[0:0] and_949_nl;
  wire[0:0] mux_731_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] and_952_nl;
  wire[0:0] mux_734_nl;
  wire[0:0] mux_733_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] and_955_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] mux_735_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] and_958_nl;
  wire[0:0] mux_740_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] and_3209_nl;
  wire[0:0] and_960_nl;
  wire[0:0] mux_743_nl;
  wire[0:0] mux_742_nl;
  wire[0:0] mux_741_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] and_962_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] mux_745_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] and_965_nl;
  wire[0:0] mux_749_nl;
  wire[0:0] mux_748_nl;
  wire[0:0] mux_747_nl;
  wire[0:0] nor_688_nl;
  wire[0:0] and_968_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] mux_751_nl;
  wire[0:0] mux_750_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] and_971_nl;
  wire[0:0] mux_755_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] mux_753_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] and_974_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_757_nl;
  wire[0:0] mux_756_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] and_977_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] mux_760_nl;
  wire[0:0] mux_759_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] and_980_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] mux_763_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] and_983_nl;
  wire[0:0] mux_767_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] and_986_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] and_989_nl;
  wire[0:0] mux_773_nl;
  wire[0:0] mux_772_nl;
  wire[0:0] mux_771_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] and_992_nl;
  wire[0:0] mux_776_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] mux_774_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] and_995_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] mux_778_nl;
  wire[0:0] mux_777_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] and_998_nl;
  wire[0:0] mux_782_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] mux_780_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] and_1001_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] mux_783_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] and_1004_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] mux_787_nl;
  wire[0:0] mux_786_nl;
  wire[0:0] and_3208_nl;
  wire[0:0] and_1006_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] and_1008_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] and_1011_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] and_1014_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] and_1017_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] and_1020_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] mux_805_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] and_1023_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] and_1026_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] mux_811_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] and_1029_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] mux_813_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] and_1032_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] and_1035_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] and_1038_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] and_1041_nl;
  wire[0:0] mux_827_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] and_1044_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] and_1047_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] and_1050_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] and_3207_nl;
  wire[0:0] and_1052_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] and_1054_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] and_1057_nl;
  wire[0:0] mux_845_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] and_1060_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] and_1063_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] and_1066_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] and_1069_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] and_1072_nl;
  wire[0:0] mux_860_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] and_1075_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] mux_861_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] and_1078_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] and_1081_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] and_1084_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] mux_871_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] and_1087_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] mux_873_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] and_1090_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] mux_877_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] and_1093_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] and_1096_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] and_1098_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] and_1100_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] and_1103_nl;
  wire[0:0] mux_893_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] and_1106_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] and_1109_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] and_1112_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] and_1115_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] and_1118_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] and_1121_nl;
  wire[0:0] mux_911_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] mux_909_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] and_1124_nl;
  wire[0:0] mux_914_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] and_1127_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] and_1130_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] and_1133_nl;
  wire[0:0] mux_923_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] and_1136_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] mux_925_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] and_1139_nl;
  wire[0:0] mux_929_nl;
  wire[0:0] mux_928_nl;
  wire[0:0] mux_927_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] and_1142_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] mux_931_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] and_3206_nl;
  wire[0:0] and_1144_nl;
  wire[0:0] mux_935_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] nor_629_nl;
  wire[0:0] and_1146_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] mux_937_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] and_1149_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] and_1152_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] mux_942_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] and_1155_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] and_1158_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] nor_624_nl;
  wire[0:0] and_1161_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] and_1164_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] and_1167_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] and_1170_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] mux_960_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] and_1173_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] and_1176_nl;
  wire[0:0] mux_968_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] mux_966_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] and_1179_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] and_1182_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] and_1185_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] and_1188_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] and_1190_nl;
  wire[0:0] mux_983_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] and_1192_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] and_1195_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] and_1198_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] and_1201_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] mux_994_nl;
  wire[0:0] mux_993_nl;
  wire[0:0] nor_609_nl;
  wire[0:0] and_1204_nl;
  wire[0:0] mux_998_nl;
  wire[0:0] mux_997_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] and_1207_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] mux_999_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] and_1210_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] and_1213_nl;
  wire[0:0] mux_1007_nl;
  wire[0:0] mux_1006_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] and_1216_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] mux_1009_nl;
  wire[0:0] mux_1008_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] and_1219_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] mux_1012_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] and_1222_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] and_1225_nl;
  wire[0:0] mux_1019_nl;
  wire[0:0] mux_1018_nl;
  wire[0:0] mux_1017_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] and_1228_nl;
  wire[0:0] mux_1022_nl;
  wire[0:0] mux_1021_nl;
  wire[0:0] mux_1020_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] and_1231_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] nor_599_nl;
  wire[0:0] and_1234_nl;
  wire[0:0] mux_1028_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] mux_1026_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] and_1236_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] mux_1030_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] and_1238_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] and_1241_nl;
  wire[0:0] mux_1037_nl;
  wire[0:0] mux_1036_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] and_1244_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] mux_1039_nl;
  wire[0:0] mux_1038_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] and_1247_nl;
  wire[0:0] mux_1043_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] mux_1041_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] and_1250_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] mux_1045_nl;
  wire[0:0] mux_1044_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] and_1253_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] mux_1047_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] and_1256_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] nor_590_nl;
  wire[0:0] and_1259_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] and_1262_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] and_1265_nl;
  wire[0:0] mux_1061_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] and_1268_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] and_1271_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] and_1274_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] and_1277_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] and_3205_nl;
  wire[0:0] and_1280_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] and_1282_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] and_1284_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] and_1287_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] and_1290_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] and_1293_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] and_1296_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] and_1299_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] and_1302_nl;
  wire[3:0] operator_8_false_3_acc_nl;
  wire[4:0] nl_operator_8_false_3_acc_nl;
  wire[1:0] LOAD_LOOP_for_if_2_for_mux_21_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_not_26_nl;
  wire[0:0] LOAD_LOOP_for_if_for_mux_4_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_mux_23_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_mux_18_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_and_200_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_or_380_nl;
  wire[1:0] LOAD_LOOP_for_if_2_for_and_198_nl;
  wire[0:0] nor_785_nl;
  wire[0:0] and_3303_nl;
  wire[0:0] and_3300_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_and_188_nl;
  wire[0:0] and_3301_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_or_176_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_and_183_nl;
  wire[0:0] nor_786_nl;
  wire[0:0] and_3299_nl;
  wire[0:0] and_3296_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_and_192_nl;
  wire[0:0] and_3297_nl;
  wire[3:0] operator_8_false_4_acc_nl;
  wire[4:0] nl_operator_8_false_4_acc_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_mux_5_nl;
  wire[9:0] LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_nl;
  wire[10:0] nl_LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_nl;
  wire[8:0] LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_1_nl;
  wire[9:0] nl_LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_1_nl;
  wire[9:0] LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_nl;
  wire[10:0] nl_LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_nl;
  wire[8:0] LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_1_nl;
  wire[9:0] nl_LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_1_nl;
  wire[4:0] operator_8_false_5_acc_nl;
  wire[5:0] nl_operator_8_false_5_acc_nl;
  wire[0:0] LOAD_LOOP_mux_1_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_mux_22_nl;
  wire[1:0] operator_8_false_1_acc_4_nl;
  wire[3:0] nl_operator_8_false_1_acc_4_nl;
  wire[2:0] operator_8_false_3_acc_2_nl;
  wire[4:0] nl_operator_8_false_3_acc_2_nl;
  wire[2:0] LOAD_LOOP_for_if_2_for_for_switch_lp_mux1h_4_nl;
  wire[1:0] operator_8_false_1_acc_3_nl;
  wire[2:0] nl_operator_8_false_1_acc_3_nl;
  wire[2:0] operator_8_false_3_operator_8_false_3_acc_nl;
  wire[3:0] nl_operator_8_false_3_operator_8_false_3_acc_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_for_switch_lp_LOAD_LOOP_for_if_2_for_for_switch_lp_and_3_nl;
  wire[0:0] LOAD_LOOP_for_if_2_for_for_switch_lp_nand_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] and_3236_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] or_180_nl;
  wire[0:0] or_177_nl;
  wire[0:0] or_192_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] and_3239_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] or_468_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] or_470_nl;
  wire[0:0] nand_33_nl;
  wire[0:0] or_469_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] or_560_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] or_559_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] or_569_nl;
  wire[0:0] nand_37_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] or_591_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] nand_279_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] or_682_nl;
  wire[0:0] or_680_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] or_731_nl;
  wire[0:0] nand_58_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] and_878_nl;
  wire[0:0] or_747_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] nand_61_nl;
  wire[0:0] nand_60_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] or_774_nl;
  wire[0:0] or_777_nl;
  wire[0:0] or_783_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] mux_504_nl;
  wire[0:0] or_782_nl;
  wire[0:0] nand_67_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] or_845_nl;
  wire[0:0] nand_79_nl;
  wire[0:0] or_872_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] nand_347_nl;
  wire[0:0] or_183_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] nand_83_nl;
  wire[0:0] or_2857_nl;
  wire[0:0] nand_81_nl;
  wire[0:0] or_899_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] or_898_nl;
  wire[0:0] nand_87_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] or_921_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] nor_695_nl;
  wire[0:0] or_928_nl;
  wire[0:0] or_935_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] or_934_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] or_447_nl;
  wire[0:0] or_446_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] or_443_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] and_840_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] nand_44_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] or_604_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] or_602_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] nand_43_nl;
  wire[0:0] or_601_nl;
  wire[0:0] nand_42_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] and_3252_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] or_189_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] and_3202_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] and_3201_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] and_3200_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] and_3199_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] and_893_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] nand_86_nl;
  wire[0:0] mux_588_nl;
  wire[0:0] or_889_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] mux_586_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] and_3222_nl;
  wire[0:0] and_3223_nl;
  wire[0:0] and_3224_nl;
  wire[8:0] LOAD_LOOP_for_if_2_for_for_if_aelse_acc_nl;
  wire[9:0] nl_LOAD_LOOP_for_if_2_for_for_if_aelse_acc_nl;
  wire[4:0] operator_8_false_6_acc_nl;
  wire[5:0] nl_operator_8_false_6_acc_nl;
  wire[0:0] nor_794_nl;
  wire[0:0] or_2906_nl;
  wire[7:0] LOAD_LOOP_for_if_2_for_for_if_index_in_mux_8_nl;
  wire[7:0] LOAD_LOOP_for_if_2_for_for_if_index_in_mux_9_nl;
  wire[7:0] LOAD_LOOP_for_if_2_for_for_if_index_in_mux_10_nl;
  wire[12:0] LOAD_LOOP_for_if_2_for_for_if_index_in_mux_11_nl;
  wire[7:0] operator_43_true_operator_43_true_acc_1_nl;
  wire[8:0] nl_operator_43_true_operator_43_true_acc_1_nl;
  wire[0:0] operator_43_true_and_1_nl;
  wire[7:0] batch_size_mux1h_14_nl;
  wire[15:0] batch_size_mux1h_15_nl;
  wire[7:0] LOAD_LOOP_for_if_for_for_index_f_mux_2_nl;
  wire[7:0] LOAD_LOOP_for_if_for_for_index_f_mux_3_nl;
  wire[7:0] pad_mux_5_nl;
  wire[13:0] pad_mux_6_nl;
  wire[7:0] LOAD_LOOP_for_mux_13_nl;
  wire[15:0] LOAD_LOOP_for_mux_14_nl;
  wire[7:0] batch_size_mux_7_nl;
  wire[15:0] batch_size_mux_8_nl;
  wire[3:0] acc_nl;
  wire[4:0] nl_acc_nl;
  wire[1:0] operator_8_false_1_mux_4_nl;
  wire[0:0] operator_8_false_1_operator_8_false_1_nor_1_nl;
  wire[0:0] operator_8_false_1_mux_5_nl;
  wire[3:0] acc_1_nl;
  wire[4:0] nl_acc_1_nl;
  wire[1:0] operator_8_false_1_mux_6_nl;
  wire[1:0] operator_8_false_1_mux_7_nl;
  wire[2:0] operator_8_false_2_mux_3_nl;
  wire[2:0] operator_8_false_3_acc_4_nl;
  wire[4:0] nl_operator_8_false_3_acc_4_nl;
  wire[1:0] operator_8_false_2_mux_4_nl;
  wire[0:0] LOAD_LOOP_for_LOAD_LOOP_for_and_2_nl;
  wire[15:0] LOAD_LOOP_for_LOAD_LOOP_for_mux_5_nl;
  wire[15:0] LOAD_LOOP_for_mux1h_9_nl;
  wire[9:0] acc_4_nl;
  wire[10:0] nl_acc_4_nl;
  wire[2:0] pad_pad_pad_nor_1_nl;
  wire[4:0] pad_mux_7_nl;
  wire[7:0] pad_mux_8_nl;
  wire[15:0] batch_size_mux1h_16_nl;
  wire[15:0] batch_size_mux1h_17_nl;
  wire[7:0] operator_8_false_3_mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_load_core_buf_linear_rsci_inst_buf_linear_rsci_oswt_unreg;
  assign nl_load_core_buf_linear_rsci_inst_buf_linear_rsci_oswt_unreg = and_dcpl_772
      & (fsm_output[2]);
  wire [4031:0] nl_load_core_buf_linear_rsci_inst_buf_linear_rsci_idat;
  assign nl_load_core_buf_linear_rsci_inst_buf_linear_rsci_idat = {buf_linear_rsci_idat_4031_4000
      , buf_linear_rsci_idat_3999_3968 , buf_linear_rsci_idat_3967_3936 , buf_linear_rsci_idat_3935_3904
      , buf_linear_rsci_idat_3903_3872 , buf_linear_rsci_idat_3871_3840 , buf_linear_rsci_idat_3839_3808
      , buf_linear_rsci_idat_3807_3776 , buf_linear_rsci_idat_3775_3744 , buf_linear_rsci_idat_3743_3712
      , buf_linear_rsci_idat_3711_3680 , buf_linear_rsci_idat_3679_3648 , buf_linear_rsci_idat_3647_3616
      , buf_linear_rsci_idat_3615_3584 , buf_linear_rsci_idat_3583_3552 , buf_linear_rsci_idat_3551_3520
      , buf_linear_rsci_idat_3519_3488 , buf_linear_rsci_idat_3487_3456 , buf_linear_rsci_idat_3455_3424
      , buf_linear_rsci_idat_3423_3392 , buf_linear_rsci_idat_3391_3360 , buf_linear_rsci_idat_3359_3328
      , buf_linear_rsci_idat_3327_3296 , buf_linear_rsci_idat_3295_3264 , buf_linear_rsci_idat_3263_3232
      , buf_linear_rsci_idat_3231_3200 , buf_linear_rsci_idat_3199_3168 , buf_linear_rsci_idat_3167_3136
      , buf_linear_rsci_idat_3135_3104 , buf_linear_rsci_idat_3103_3072 , buf_linear_rsci_idat_3071_3040
      , buf_linear_rsci_idat_3039_3008 , buf_linear_rsci_idat_3007_2976 , buf_linear_rsci_idat_2975_2944
      , buf_linear_rsci_idat_2943_2912 , buf_linear_rsci_idat_2911_2880 , buf_linear_rsci_idat_2879_2848
      , buf_linear_rsci_idat_2847_2816 , buf_linear_rsci_idat_2815_2784 , buf_linear_rsci_idat_2783_2752
      , buf_linear_rsci_idat_2751_2720 , buf_linear_rsci_idat_2719_2688 , buf_linear_rsci_idat_2687_2656
      , buf_linear_rsci_idat_2655_2624 , buf_linear_rsci_idat_2623_2592 , buf_linear_rsci_idat_2591_2560
      , buf_linear_rsci_idat_2559_2528 , buf_linear_rsci_idat_2527_2496 , buf_linear_rsci_idat_2495_2464
      , buf_linear_rsci_idat_2463_2432 , buf_linear_rsci_idat_2431_2400 , buf_linear_rsci_idat_2399_2368
      , buf_linear_rsci_idat_2367_2336 , buf_linear_rsci_idat_2335_2304 , buf_linear_rsci_idat_2303_2272
      , buf_linear_rsci_idat_2271_2240 , buf_linear_rsci_idat_2239_2208 , buf_linear_rsci_idat_2207_2176
      , buf_linear_rsci_idat_2175_2144 , buf_linear_rsci_idat_2143_2112 , buf_linear_rsci_idat_2111_2080
      , buf_linear_rsci_idat_2079_2048 , buf_linear_rsci_idat_2047_2016 , buf_linear_rsci_idat_2015_1984
      , buf_linear_rsci_idat_1983_1952 , buf_linear_rsci_idat_1951_1920 , buf_linear_rsci_idat_1919_1888
      , buf_linear_rsci_idat_1887_1856 , buf_linear_rsci_idat_1855_1824 , buf_linear_rsci_idat_1823_1792
      , buf_linear_rsci_idat_1791_1760 , buf_linear_rsci_idat_1759_1728 , buf_linear_rsci_idat_1727_1696
      , buf_linear_rsci_idat_1695_1664 , buf_linear_rsci_idat_1663_1632 , buf_linear_rsci_idat_1631_1600
      , buf_linear_rsci_idat_1599_1568 , buf_linear_rsci_idat_1567_1536 , buf_linear_rsci_idat_1535_1504
      , buf_linear_rsci_idat_1503_1472 , buf_linear_rsci_idat_1471_1440 , buf_linear_rsci_idat_1439_1408
      , buf_linear_rsci_idat_1407_1376 , buf_linear_rsci_idat_1375_1344 , buf_linear_rsci_idat_1343_1312
      , buf_linear_rsci_idat_1311_1280 , buf_linear_rsci_idat_1279_1248 , buf_linear_rsci_idat_1247_1216
      , buf_linear_rsci_idat_1215_1184 , buf_linear_rsci_idat_1183_1152 , buf_linear_rsci_idat_1151_1120
      , buf_linear_rsci_idat_1119_1088 , buf_linear_rsci_idat_1087_1056 , buf_linear_rsci_idat_1055_1024
      , buf_linear_rsci_idat_1023_992 , buf_linear_rsci_idat_991_960 , buf_linear_rsci_idat_959_928
      , buf_linear_rsci_idat_927_896 , buf_linear_rsci_idat_895_864 , buf_linear_rsci_idat_863_832
      , buf_linear_rsci_idat_831_800 , buf_linear_rsci_idat_799_768 , buf_linear_rsci_idat_767_736
      , buf_linear_rsci_idat_735_704 , buf_linear_rsci_idat_703_672 , buf_linear_rsci_idat_671_640
      , buf_linear_rsci_idat_639_608 , buf_linear_rsci_idat_607_576 , buf_linear_rsci_idat_575_544
      , buf_linear_rsci_idat_543_512 , buf_linear_rsci_idat_511_480 , buf_linear_rsci_idat_479_448
      , buf_linear_rsci_idat_447_416 , buf_linear_rsci_idat_415_384 , buf_linear_rsci_idat_383_352
      , buf_linear_rsci_idat_351_320 , buf_linear_rsci_idat_319_288 , buf_linear_rsci_idat_287_256
      , buf_linear_rsci_idat_255_224 , buf_linear_rsci_idat_223_192 , buf_linear_rsci_idat_191_160
      , buf_linear_rsci_idat_159_128 , buf_linear_rsci_idat_127_96 , buf_linear_rsci_idat_95_64
      , buf_linear_rsci_idat_63_32 , buf_linear_rsci_idat_31_0};
  wire [0:0] nl_load_core_plm_kernel_rsci_inst_plm_kernel_rsci_oswt_unreg;
  assign nl_load_core_plm_kernel_rsci_inst_plm_kernel_rsci_oswt_unreg = or_tmp_4
      & and_dcpl_764 & (fsm_output[2]);
  wire [1567:0] nl_load_core_plm_kernel_rsci_inst_plm_kernel_rsci_idat;
  assign nl_load_core_plm_kernel_rsci_inst_plm_kernel_rsci_idat = {plm_kernel_rsci_idat_1567_1536
      , plm_kernel_rsci_idat_1535_1504 , plm_kernel_rsci_idat_1503_1472 , plm_kernel_rsci_idat_1471_1440
      , plm_kernel_rsci_idat_1439_1408 , plm_kernel_rsci_idat_1407_1376 , plm_kernel_rsci_idat_1375_1344
      , plm_kernel_rsci_idat_1343_1312 , plm_kernel_rsci_idat_1311_1280 , plm_kernel_rsci_idat_1279_1248
      , plm_kernel_rsci_idat_1247_1216 , plm_kernel_rsci_idat_1215_1184 , plm_kernel_rsci_idat_1183_1152
      , plm_kernel_rsci_idat_1151_1120 , plm_kernel_rsci_idat_1119_1088 , plm_kernel_rsci_idat_1087_1056
      , plm_kernel_rsci_idat_1055_1024 , plm_kernel_rsci_idat_1023_992 , plm_kernel_rsci_idat_991_960
      , plm_kernel_rsci_idat_959_928 , plm_kernel_rsci_idat_927_896 , plm_kernel_rsci_idat_895_864
      , plm_kernel_rsci_idat_863_832 , plm_kernel_rsci_idat_831_800 , plm_kernel_rsci_idat_799_768
      , plm_kernel_rsci_idat_767_736 , plm_kernel_rsci_idat_735_704 , plm_kernel_rsci_idat_703_672
      , plm_kernel_rsci_idat_671_640 , plm_kernel_rsci_idat_639_608 , plm_kernel_rsci_idat_607_576
      , plm_kernel_rsci_idat_575_544 , plm_kernel_rsci_idat_543_512 , plm_kernel_rsci_idat_511_480
      , plm_kernel_rsci_idat_479_448 , plm_kernel_rsci_idat_447_416 , plm_kernel_rsci_idat_415_384
      , plm_kernel_rsci_idat_383_352 , plm_kernel_rsci_idat_351_320 , plm_kernel_rsci_idat_319_288
      , plm_kernel_rsci_idat_287_256 , plm_kernel_rsci_idat_255_224 , plm_kernel_rsci_idat_223_192
      , plm_kernel_rsci_idat_191_160 , plm_kernel_rsci_idat_159_128 , plm_kernel_rsci_idat_127_96
      , plm_kernel_rsci_idat_95_64 , plm_kernel_rsci_idat_63_32 , plm_kernel_rsci_idat_31_0};
  wire [0:0] nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_oswt_unreg;
  assign nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_oswt_unreg = (~((~(LOAD_LOOP_for_asn_2_itm_1
      & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]))) & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1])))
      & LOAD_BATCH_LOOP_and_3_tmp & (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2)
      & (fsm_output[2]);
  wire [66:0] nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat;
  assign nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat = {19'b0110000000000000000
      , dma_read_ctrl_rsci_idat_47_32 , 16'b0000000000000000 , dma_read_ctrl_rsci_idat_15_0};
  wire[0:0] mux_298_nl;
  wire[0:0] mux_297_nl;
  wire [0:0] nl_load_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg;
  assign mux_297_nl = MUX_s_1_2_2((~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1])),
      (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]), lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2);
  assign mux_298_nl = MUX_s_1_2_2(or_dcpl_34, mux_297_nl, and_3198_cse);
  assign nl_load_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg = (~
      mux_298_nl) & and_dcpl_738 & (fsm_output[2]);
  wire [0:0] nl_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_inst_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg;
  assign nl_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_inst_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg
      = or_tmp_4 & and_dcpl_182 & LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt & LOAD_LOOP_for_if_2_for_for_asn_itm_2
      & LOAD_BATCH_LOOP_stage_0_3 & (fsm_output[2]);
  wire [0:0] nl_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_inst_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1;
  assign nl_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_inst_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1
      = or_tmp_4 & and_dcpl_176 & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]))
      & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2 & (~ LOAD_LOOP_for_if_2_for_for_asn_itm_2)
      & LOAD_BATCH_LOOP_stage_0_3 & (fsm_output[2]);
  esp_acc_conv2dlb_cxx_catapult_load_core_conf_info_rsci load_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt(reg_conf_info_rsci_irdy_core_psct_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_buf_linear_rsci load_core_buf_linear_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .buf_linear_rsc_dat(buf_linear_rsc_dat),
      .buf_linear_rsc_vld(buf_linear_rsc_vld),
      .buf_linear_rsc_rdy(buf_linear_rsc_rdy),
      .core_wen(core_wen),
      .buf_linear_rsci_oswt_unreg(nl_load_core_buf_linear_rsci_inst_buf_linear_rsci_oswt_unreg[0:0]),
      .buf_linear_rsci_bawt(buf_linear_rsci_bawt),
      .buf_linear_rsci_iswt0(reg_buf_linear_rsci_ivld_core_psct_cse),
      .buf_linear_rsci_wen_comp(buf_linear_rsci_wen_comp),
      .buf_linear_rsci_idat(nl_load_core_buf_linear_rsci_inst_buf_linear_rsci_idat[4031:0])
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_plm_kernel_rsci load_core_plm_kernel_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_kernel_rsc_dat(plm_kernel_rsc_dat),
      .plm_kernel_rsc_vld(plm_kernel_rsc_vld),
      .plm_kernel_rsc_rdy(plm_kernel_rsc_rdy),
      .core_wen(core_wen),
      .plm_kernel_rsci_oswt_unreg(nl_load_core_plm_kernel_rsci_inst_plm_kernel_rsci_oswt_unreg[0:0]),
      .plm_kernel_rsci_bawt(plm_kernel_rsci_bawt),
      .plm_kernel_rsci_iswt0(reg_plm_kernel_rsci_ivld_core_psct_cse),
      .plm_kernel_rsci_wen_comp(plm_kernel_rsci_wen_comp),
      .plm_kernel_rsci_idat(nl_load_core_plm_kernel_rsci_inst_plm_kernel_rsci_idat[1567:0])
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_ctrl_rsci load_core_dma_read_ctrl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dma_read_ctrl_rsci_oswt_unreg(nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_oswt_unreg[0:0]),
      .dma_read_ctrl_rsci_bawt(dma_read_ctrl_rsci_bawt),
      .dma_read_ctrl_rsci_iswt0(reg_dma_read_ctrl_rsci_ivld_core_psct_cse),
      .dma_read_ctrl_rsci_irdy_mxwt(dma_read_ctrl_rsci_irdy_mxwt),
      .dma_read_ctrl_rsci_idat(nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat[66:0])
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_dma_read_chnl_rsci load_core_dma_read_chnl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .core_wen(core_wen),
      .dma_read_chnl_rsci_oswt_unreg(nl_load_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg[0:0]),
      .dma_read_chnl_rsci_bawt(dma_read_chnl_rsci_bawt),
      .dma_read_chnl_rsci_iswt0(reg_dma_read_chnl_rsci_irdy_core_psct_cse),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .dma_read_chnl_rsci_idat_mxwt(dma_read_chnl_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_done_rsci load_core_done_rsci_inst (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt(reg_done_rsci_ivld_core_psct_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1
      load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_inst (
      .clk(clk),
      .rst(rst),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg(nl_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_inst_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg[0:0]),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0(reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1(nl_load_core_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_1_inst_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_oswt_unreg_1[0:0]),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1(reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_iff),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_pff(and_2372_rmff),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_iswt0_1_pff(and_2370_rmff)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_staller load_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .buf_linear_rsci_wen_comp(buf_linear_rsci_wen_comp),
      .plm_kernel_rsci_wen_comp(plm_kernel_rsci_wen_comp),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core_core_fsm load_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output),
      .LOAD_BATCH_LOOP_C_0_tr0(and_dcpl_24)
    );
  assign or_1869_nl = LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (~ (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0]));
  assign mux_1098_nl = MUX_s_1_2_2(or_1869_nl, exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2,
      or_75_cse);
  assign and_1304_tmp = (~ mux_1098_nl) & and_3266_cse;
  assign and_2370_rmff = and_dcpl_739 & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2
      & (~ LOAD_LOOP_for_if_2_for_for_asn_itm_1) & (fsm_output[2]);
  assign and_2372_rmff = and_dcpl_739 & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2
      & LOAD_LOOP_for_if_2_for_for_asn_itm_1 & (fsm_output[2]);
  assign and_808_nl = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 & mux_tmp_260;
  assign mux_279_nl = MUX_s_1_2_2(and_808_nl, and_tmp_22, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]);
  assign mux_1159_itm = MUX_s_1_2_2(or_tmp_340, mux_279_nl, nor_113_cse);
  assign and_3198_cse = LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st_1 & LOAD_LOOP_for_if_2_for_for_asn_itm_1;
  assign LOAD_LOOP_for_if_2_for_for_if_index_in_mux_rmff = MUX_v_14_2_2(LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d_reg, or_tmp_2041);
  assign or_2436_nl = (~ (fsm_output[2])) | or_dcpl_129 | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2)
      | LOAD_LOOP_for_if_2_for_for_asn_itm_1;
  assign LOAD_LOOP_for_if_2_for_for_else_index_in_mux_rmff = MUX_v_14_2_2(LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d_reg, or_2436_nl);
  assign LOAD_LOOP_for_if_2_for_for_if_mux_rmff = MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_mx0w0,
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d_reg, or_tmp_2041);
  assign or_2860_cse = (~((~ LOAD_LOOP_for_if_3_equal_tmp) | (operator_8_false_6_acc_tmp[8:5]!=4'b0000)))
      | (LOAD_LOOP_for_acc_2_tmp[5]);
  assign or_513_cse = (~((operator_8_false_7_acc_tmp[8:5]!=4'b0000) | (~ LOAD_LOOP_if_equal_tmp)))
      | (LOAD_LOOP_acc_tmp[5]);
  assign LOAD_LOOP_for_if_for_and_cse = core_wen & (fsm_output[2]) & LOAD_BATCH_LOOP_and_3_tmp;
  assign LOAD_LOOP_for_if_2_for_if_and_128_cse = core_wen & (~((~ (fsm_output[2]))
      | or_dcpl_135));
  assign and_3197_cse = ((~ LOAD_LOOP_for_if_for_for_if_equal_tmp) | (operator_8_false_1_acc_tmp[8:3]!=6'b000000))
      & operator_8_false_4_acc_itm_3_1;
  assign or_539_cse = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b10)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign mux_333_nl = MUX_s_1_2_2(or_750_cse, (~ or_750_cse), dma_read_ctrl_rsci_irdy_mxwt);
  assign mux_335_cse = MUX_s_1_2_2((~ or_750_cse), mux_333_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign and_834_cse = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 & mux_335_cse;
  assign LOAD_LOOP_for_if_2_for_and_205_cse = core_wen & (~((~ (fsm_output[2])) |
      mux_tmp_353 | or_dcpl_146));
  assign LOAD_LOOP_for_if_for_and_2_cse = core_wen & (fsm_output[2]) & LOAD_BATCH_LOOP_and_4_tmp;
  assign nor_752_cse = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0!=2'b11));
  assign or_631_cse = (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00);
  assign or_632_cse = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00);
  assign and_849_nl = or_634_cse & mux_tmp_399;
  assign mux_401_nl = MUX_s_1_2_2(mux_tmp_399, and_849_nl, nor_tmp_172);
  assign LOAD_LOOP_for_if_for_and_3_cse = core_wen & (fsm_output[2]) & mux_401_nl
      & LOAD_BATCH_LOOP_and_4_tmp;
  assign LOAD_LOOP_for_if_2_for_for_col_and_2_cse = core_wen & and_3158_cse;
  assign or_654_cse = buf_linear_rsci_bawt | (~ LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3)
      | (~ exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0[1])
      | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0[0]);
  assign nor_178_cse = ~(LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (~ (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0])));
  assign and_3195_cse = or_tmp_154 & (~ LOAD_LOOP_for_if_2_for_equal_tmp_2_1) & (LOAD_LOOP_for_if_2_for_mux1h_378_tmp==2'b11);
  assign LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse = (LOAD_BATCH_LOOP_acc_tmp[4])
      | LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_nor_tmp;
  assign or_750_cse = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0!=2'b11)
      | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2;
  assign or_755_cse = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign and_3192_cse = (~ LOAD_LOOP_for_asn_6_itm_1) & LOAD_LOOP_for_if_2_for_equal_tmp_1_1;
  assign nor_225_cse = ~(nor_tmp_50 | (~ LOAD_LOOP_for_if_2_for_equal_tmp_1_1));
  assign LOAD_LOOP_for_if_for_for_and_111_cse = core_wen & (~((~ (fsm_output[2]))
      | or_dcpl_128 | or_dcpl_34));
  assign LOAD_LOOP_for_and_2_cse = core_wen & (fsm_output[2]);
  assign or_766_nl = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b11)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign nand_64_nl = ~(LOAD_LOOP_for_if_2_for_and_195_ssc_1 & (~ and_834_cse));
  assign mux_480_nl = MUX_s_1_2_2(nand_64_nl, and_834_cse, and_3195_cse);
  assign mux_481_cse = MUX_s_1_2_2(or_766_nl, mux_480_nl, nor_37_cse);
  assign LOAD_LOOP_for_if_2_for_for_and_257_cse = core_wen & (~((~ (fsm_output[2]))
      | mux_tmp_353 | or_dcpl_136));
  assign nor_566_cse = ~(buf_linear_rsci_bawt | (~ LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3)
      | (~ exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0[1])
      | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0[0]));
  assign mux_491_cse = MUX_s_1_2_2(mux_tmp_486, mux_tmp_484, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_497_cse = MUX_s_1_2_2(nand_tmp_66, nand_tmp_65, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_510_cse = MUX_s_1_2_2(mux_tmp_505, mux_tmp_502, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign or_771_cse = nor_566_cse | LOAD_BATCH_LOOP_stage_0_3;
  assign or_810_cse = (~ operator_8_false_5_acc_itm_4_1) | LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_1_LOAD_LOOP_for_if_2_for_if_1_nor_tmp;
  assign LOAD_LOOP_for_if_2_for_for_and_259_cse = core_wen & (~((~ (fsm_output[2]))
      | (~ or_tmp_4) | or_dcpl_122 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1])
      | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2) | and_dcpl_186 | (~
      LOAD_BATCH_LOOP_stage_0_3)));
  assign operator_8_false_and_cse = core_wen & (or_tmp_2314 | or_tmp_2315);
  assign LOAD_LOOP_for_if_2_for_if_and_132_cse = core_wen & LOAD_BATCH_LOOP_and_3_tmp;
  assign LOAD_LOOP_for_if_for_for_n_and_1_cse = core_wen & ((fsm_output[1]) | or_tmp_2337);
  assign or_75_cse = (~ LOAD_BATCH_LOOP_and_3_tmp) | LOAD_BATCH_LOOP_asn_itm_1;
  assign nor_32_cse = ~(LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_1_LOAD_LOOP_for_if_2_for_if_1_nor_tmp
      | (~ operator_8_false_5_acc_itm_4_1));
  assign and_cse = core_wen & (~ (fsm_output[2]));
  assign LOAD_LOOP_fl_and_cse = core_wen & ((fsm_output[1]) | or_tmp_2354);
  assign mux_609_cse = MUX_s_1_2_2(mux_tmp_604, nor_tmp_291, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_606_nl = MUX_s_1_2_2(mux_tmp_604, nor_tmp_291, nor_tmp_54);
  assign mux_608_nl = MUX_s_1_2_2(mux_609_cse, mux_606_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_610_nl = MUX_s_1_2_2(mux_609_cse, mux_608_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_611_nl = MUX_s_1_2_2(mux_609_cse, mux_610_nl, nor_752_cse);
  assign LOAD_LOOP_for_and_5_cse = core_wen & (~((~ mux_611_nl) & and_3266_cse))
      & LOAD_BATCH_LOOP_and_4_tmp;
  assign LOAD_LOOP_for_and_9_cse = core_wen & ((fsm_output[1]) | or_tmp_2314) & (exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0
      | (~ or_tmp_2314));
  assign or_1873_tmp = mux_tmp_353 | and_dcpl_779 | (~ lfst_exit_LOAD_LOOP_for_1_lpi_2)
      | and_dcpl_778 | (~ lfst_exit_LOAD_LOOP_sva);
  assign mux_619_cse = MUX_s_1_2_2(mux_tmp_614, mux_tmp_612, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign and_3158_cse = LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign or_941_cse = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0!=2'b10);
  assign or_939_cse = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]!=3'b000);
  assign and_3220_cse = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]==3'b111);
  assign or_950_cse = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]!=3'b001);
  assign nor_302_cse = ~((LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]!=3'b110));
  assign nor_304_cse = ~((LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]!=3'b010));
  assign or_960_cse = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]!=3'b101);
  assign nor_307_cse = ~((LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]!=3'b011));
  assign or_967_cse = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2:0]!=3'b100);
  assign nand_225_cse = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 & or_tmp_4);
  assign nand_224_cse = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 & or_tmp_4);
  assign nand_222_cse = ~(or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b10));
  assign nand_223_cse = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 & or_tmp_4);
  assign nand_218_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 & or_tmp_4);
  assign nand_215_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 & or_tmp_4);
  assign nand_213_cse = ~(or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])));
  assign nand_214_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 & or_tmp_4);
  assign nand_212_cse = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      & or_tmp_4);
  assign nand_199_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 & or_tmp_4);
  assign nand_197_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 & or_tmp_4);
  assign nand_195_cse = ~(or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b110));
  assign nand_196_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 & or_tmp_4);
  assign nand_194_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      & or_tmp_4);
  assign nand_167_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 & or_tmp_4);
  assign nand_165_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 & or_tmp_4);
  assign nand_164_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 & or_tmp_4);
  assign nand_163_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      & or_tmp_4);
  assign or_481_cse = (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b10);
  assign nl_operator_8_false_3_acc_nl = ({1'b1 , LOAD_LOOP_for_if_for_m_2_0_sva_1_mx0w1})
      + 4'b0001;
  assign operator_8_false_3_acc_nl = nl_operator_8_false_3_acc_nl[3:0];
  assign exit_LOAD_LOOP_for_if_for_lpi_2_dfm_mx0w0 = (~ (readslicef_4_1_3(operator_8_false_3_acc_nl)))
      | exit_LOAD_LOOP_for_if_for_sva_1_mx0w0;
  assign exit_LOAD_LOOP_lpi_2_dfm_1_mx0w0 = (LOAD_LOOP_acc_tmp[5]) | exit_LOAD_LOOP_sva_3;
  assign LOAD_LOOP_for_if_2_for_equal_tmp_2_mx0w0 = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1
      & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1==2'b00);
  assign LOAD_LOOP_for_if_2_for_mux_21_nl = MUX_v_2_2_2(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0_mx0w0,
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0, or_75_cse);
  assign LOAD_LOOP_for_if_2_for_not_26_nl = ~ exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1;
  assign lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1 = MUX_v_2_2_2(2'b00,
      LOAD_LOOP_for_if_2_for_mux_21_nl, LOAD_LOOP_for_if_2_for_not_26_nl);
  assign LOAD_LOOP_for_if_for_mux_4_nl = MUX_s_1_2_2(exit_LOAD_LOOP_for_if_for_lpi_2_dfm_mx0w0,
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm, and_3197_cse);
  assign exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0 = LOAD_LOOP_for_if_for_mux_4_nl
      & exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_mx0w0;
  assign LOAD_LOOP_for_if_2_for_equal_tmp_mx0w0 = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1[1])
      & (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1[0])));
  assign LOAD_LOOP_for_if_2_for_equal_tmp_1_mx0w0 = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1==2'b11)
      & (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1);
  assign LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_if_1_LOAD_LOOP_for_if_2_for_for_if_1_nor_tmp
      = ~((~((LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1 == (operator_8_false_4_acc_psp_sva_1[4:0]))
      & (operator_8_false_4_acc_psp_sva_1[7:5]==3'b000))) | (operator_8_false_4_acc_psp_sva_1[8]));
  assign nl_LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1 = LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1
      + 5'b00001;
  assign LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1 = nl_LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1[4:0];
  assign exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0 = (~ operator_8_false_6_acc_itm_4_1)
      | LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_if_1_LOAD_LOOP_for_if_2_for_for_if_1_nor_tmp;
  assign nl_LOAD_LOOP_for_if_2_for_row_4_0_sva_1_mx0w1 = LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1
      + 5'b00001;
  assign LOAD_LOOP_for_if_2_for_row_4_0_sva_1_mx0w1 = nl_LOAD_LOOP_for_if_2_for_row_4_0_sva_1_mx0w1[4:0];
  assign LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_1_LOAD_LOOP_for_if_2_for_if_1_nor_tmp
      = ~((~((LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1 == (operator_8_false_5_acc_psp_sva_1[4:0]))
      & (operator_8_false_5_acc_psp_sva_1[7:5]==3'b000))) | (operator_8_false_5_acc_psp_sva_1[8]));
  assign nl_LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1 = LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_mx1
      + 3'b001;
  assign LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1 = nl_LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1[2:0];
  assign LOAD_LOOP_for_if_for_for_if_equal_tmp = LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_mx1
      == (operator_8_false_1_acc_tmp[2:0]);
  assign exit_LOAD_LOOP_for_if_for_for_sva_mx0w0 = ~((~(LOAD_LOOP_for_if_for_for_if_equal_tmp
      & LOAD_LOOP_for_if_for_for_if_nor_cse_sva_1)) | (operator_8_false_1_acc_tmp[8]));
  assign exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_mx0w0 = (~ operator_8_false_4_acc_itm_3_1)
      | exit_LOAD_LOOP_for_if_for_for_sva_mx0w0;
  assign nl_LOAD_LOOP_for_if_for_m_2_0_sva_1_mx0w1 = LOAD_LOOP_for_if_for_m_2_0_lpi_2_mx1
      + 3'b001;
  assign LOAD_LOOP_for_if_for_m_2_0_sva_1_mx0w1 = nl_LOAD_LOOP_for_if_for_m_2_0_sva_1_mx0w1[2:0];
  assign exit_LOAD_LOOP_for_if_for_sva_1_mx0w0 = ~((~((LOAD_LOOP_for_if_for_m_2_0_lpi_2_mx1
      == (operator_8_false_1_acc_tmp[2:0])) & LOAD_LOOP_for_if_for_for_if_nor_cse_sva_1))
      | (operator_8_false_1_acc_tmp[8]));
  assign LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_mx0w0 = (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1
      == LOAD_LOOP_for_print_buf_lpi_2_mx1_4_0) & (LOAD_LOOP_for_print_buf_lpi_2_mx2_7_5==3'b000);
  assign LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_mx0w1 = LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_itm_9_1
      & LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_itm_9_1 & (~(LOAD_LOOP_for_if_2_for_for_if_aelse_acc_itm_8
      | (z_out_11[8])));
  assign LOAD_LOOP_for_if_2_for_mux_23_nl = MUX_s_1_2_2(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2_mx0w0,
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2, or_75_cse);
  assign lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1 = LOAD_LOOP_for_if_2_for_mux_23_nl
      & (~ exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1);
  assign nl_LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3_mx0w0
      = conv_u2u_1_3(LOAD_LOOP_for_if_2_for_for_acc_2_psp_1[3]) + LOAD_LOOP_for_if_2_for_for_row_norm_2_0_lpi_2_dfm_1;
  assign LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3_mx0w0
      = nl_LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3_mx0w0[2:0];
  assign exit_LOAD_LOOP_for_lpi_2_dfm_3_mx0w0 = ((LOAD_LOOP_for_acc_2_tmp[5]) | (~((~(LOAD_LOOP_for_if_3_equal_tmp
      & (operator_8_false_6_acc_tmp[7:5]==3'b000))) | (operator_8_false_6_acc_tmp[8]))))
      & exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_3 & LOAD_LOOP_for_if_2_for_equal_tmp_2_mx0w0;
  assign exitL_exit_LOAD_LOOP_for_if_2_for_sva_1_mx0w0 = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2_mx0w0
      | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0_mx0w0!=2'b00));
  assign LOAD_LOOP_for_if_2_for_mux_18_nl = MUX_s_1_2_2(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2,
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2_mx0w0 = (LOAD_LOOP_for_if_2_for_mux_18_nl
      & (~(LOAD_LOOP_for_if_2_for_or_tmp_1 | LOAD_LOOP_for_if_2_for_and_195_ssc_1)))
      | LOAD_LOOP_for_if_2_for_and_181_cse_1;
  assign LOAD_LOOP_for_if_2_for_and_199_cse = (~ dma_read_ctrl_rsci_irdy_mxwt) &
      LOAD_LOOP_for_if_2_for_or_tmp_1;
  assign LOAD_LOOP_for_if_2_for_and_200_nl = dma_read_ctrl_rsci_irdy_mxwt & LOAD_LOOP_for_if_2_for_or_tmp_1;
  assign LOAD_LOOP_for_if_2_for_or_380_nl = ((~ exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_1)
      & LOAD_LOOP_for_if_2_for_equal_tmp_1) | LOAD_LOOP_for_if_2_for_and_180_cse_1
      | LOAD_LOOP_for_if_2_for_nor_tmp_1;
  assign LOAD_LOOP_for_if_2_for_mux1h_378_tmp = MUX1HOT_v_2_3_2(2'b01, 2'b10, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_1_0,
      {LOAD_LOOP_for_if_2_for_and_199_cse , LOAD_LOOP_for_if_2_for_and_200_nl , LOAD_LOOP_for_if_2_for_or_380_nl});
  assign LOAD_LOOP_for_if_2_for_and_198_nl = LOAD_LOOP_for_if_2_for_mux1h_378_tmp
      & (signext_2_1(~ LOAD_LOOP_for_if_2_for_equal_tmp_2_1)) & (signext_2_1(~ LOAD_LOOP_for_if_2_for_and_181_cse_1));
  assign lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0_mx0w0 = MUX_v_2_2_2(LOAD_LOOP_for_if_2_for_and_198_nl,
      2'b11, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign or_2893_tmp = or_dcpl_395 | ((~ LOAD_LOOP_for_if_for_for_and_tmp_1) & LOAD_LOOP_for_if_2_for_equal_tmp_1)
      | LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
  assign LOAD_LOOP_for_if_2_for_and_187_tmp = LOAD_LOOP_for_if_for_for_and_tmp_1
      & LOAD_LOOP_for_if_2_for_equal_tmp_1;
  assign nor_785_nl = ~(LOAD_LOOP_for_if_2_for_and_187_tmp | or_2893_tmp);
  assign and_3303_nl = LOAD_LOOP_for_if_2_for_and_187_tmp & (~ or_2893_tmp);
  assign LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3_mx0w0 = MUX1HOT_v_3_3_2((signext_3_1(~
      dma_read_ctrl_rsci_irdy_mxwt)), LOAD_LOOP_for_if_for_m_2_0_sva_1_1, LOAD_LOOP_for_if_for_m_2_0_lpi_2,
      {nor_785_nl , and_3303_nl , or_2893_tmp});
  assign or_2895_tmp = or_dcpl_395 | (exit_LOAD_LOOP_for_if_for_for_sva_1 & LOAD_LOOP_for_if_2_for_and_176_m1c_1)
      | LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
  assign and_3300_nl = LOAD_LOOP_for_if_2_for_or_tmp_1 & (~ or_2895_tmp);
  assign LOAD_LOOP_for_if_2_for_and_188_nl = LOAD_LOOP_for_if_2_for_and_176_m1c_1
      & (~ or_2895_tmp);
  assign and_3301_nl = exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_1 & LOAD_LOOP_for_if_2_for_equal_tmp_1
      & (~ or_2895_tmp);
  assign LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4_mx0w0 = MUX1HOT_v_3_4_2((signext_3_1(~
      dma_read_ctrl_rsci_irdy_mxwt)), LOAD_LOOP_for_if_for_for_n_2_0_sva_1_1, LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_2_1,
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2, {and_3300_nl , LOAD_LOOP_for_if_2_for_and_188_nl
      , and_3301_nl , or_2895_tmp});
  assign sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1_mx0w0 = LOAD_LOOP_for_if_2_for_mux_11_itm_1
      & (~ LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign LOAD_LOOP_for_if_2_for_or_176_nl = LOAD_LOOP_for_if_2_for_or_tmp_1 | LOAD_LOOP_for_if_2_for_equal_tmp_1
      | LOAD_LOOP_for_if_2_for_nor_tmp_1 | LOAD_LOOP_for_if_2_for_and_180_cse_1 |
      ((~ LOAD_LOOP_for_if_2_for_for_and_250_tmp_1) & LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign LOAD_LOOP_for_if_2_for_and_183_nl = LOAD_LOOP_for_if_2_for_for_and_250_tmp_1
      & LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
  assign LOAD_LOOP_for_print_buf_lpi_2_dfm_3_mx0w0 = MUX1HOT_v_8_3_2(LOAD_LOOP_for_print_buf_lpi_2,
      (z_out_13[7:0]), LOAD_LOOP_for_print_buf_sva_1_1, {LOAD_LOOP_for_if_2_for_or_176_nl
      , LOAD_LOOP_for_if_2_for_and_181_cse_1 , LOAD_LOOP_for_if_2_for_and_183_nl});
  assign or_2899_tmp = or_dcpl_401 | (LOAD_LOOP_for_if_2_for_equal_tmp_2_1 & (~ LOAD_LOOP_for_if_2_for_for_and_251_tmp_1))
      | LOAD_LOOP_for_if_2_for_equal_tmp_1;
  assign LOAD_LOOP_for_if_2_for_and_191_tmp = LOAD_LOOP_for_if_2_for_for_and_251_tmp_1
      & LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
  assign nor_786_nl = ~(LOAD_LOOP_for_if_2_for_and_191_tmp | or_2899_tmp);
  assign and_3299_nl = LOAD_LOOP_for_if_2_for_and_191_tmp & (~ or_2899_tmp);
  assign LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3_mx0w0 = MUX1HOT_v_5_3_2((signext_5_1(~
      exitL_exit_LOAD_CTRL_LOOP2_lpi_2_dfm_1)), LOAD_LOOP_for_if_2_for_row_4_0_sva_1_1,
      LOAD_LOOP_for_if_2_for_row_4_0_lpi_2, {nor_786_nl , and_3299_nl , or_2899_tmp});
  assign or_2901_tmp = or_dcpl_401 | (exit_LOAD_LOOP_for_if_2_for_for_sva_1 & LOAD_LOOP_for_if_2_for_and_178_m1c_1)
      | LOAD_LOOP_for_if_2_for_equal_tmp_1;
  assign and_3296_nl = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 & (~ or_2901_tmp);
  assign LOAD_LOOP_for_if_2_for_and_192_nl = LOAD_LOOP_for_if_2_for_and_178_m1c_1
      & (~ or_2901_tmp);
  assign and_3297_nl = exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_1 & LOAD_LOOP_for_if_2_for_equal_tmp_2_1
      & (~ or_2901_tmp);
  assign LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4_mx0w0 = MUX1HOT_v_5_4_2((signext_5_1(~
      exitL_exit_LOAD_CTRL_LOOP2_lpi_2_dfm_1)), LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_1,
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_2_1, LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2,
      {and_3296_nl , LOAD_LOOP_for_if_2_for_and_192_nl , and_3297_nl , or_2901_tmp});
  assign LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_mx1 = MUX_v_3_2_2(LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4_mx0w0,
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2, or_75_cse);
  assign LOAD_LOOP_for_if_for_m_2_0_lpi_2_mx1 = MUX_v_3_2_2(LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3_mx0w0,
      LOAD_LOOP_for_if_for_m_2_0_lpi_2, or_75_cse);
  assign LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1 = MUX_v_5_2_2(LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4_mx0w0,
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2, or_75_cse);
  assign LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1 = MUX_v_5_2_2(LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3_mx0w0,
      LOAD_LOOP_for_if_2_for_row_4_0_lpi_2, or_75_cse);
  assign sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_mx1 = MUX_s_1_2_2(sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1_mx0w0,
      sfi_operator_8_false_operator_8_false_nor_cse_lpi_2, or_75_cse);
  assign LOAD_LOOP_for_print_buf_lpi_2_mx1_4_0 = MUX_v_5_2_2((LOAD_LOOP_for_print_buf_lpi_2_dfm_3_mx0w0[4:0]),
      (LOAD_LOOP_for_print_buf_lpi_2[4:0]), or_75_cse);
  assign LOAD_LOOP_for_print_buf_lpi_2_mx2_7_5 = MUX_v_3_2_2((LOAD_LOOP_for_print_buf_lpi_2_dfm_3_mx0w0[7:5]),
      (LOAD_LOOP_for_print_buf_lpi_2[7:5]), or_75_cse);
  assign lfst_exit_LOAD_LOOP_sva_dfm_1_mx0w1 = (LOAD_BATCH_LOOP_acc_tmp[4]) | LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_nor_tmp
      | (~ exit_LOAD_LOOP_lpi_2_dfm_4);
  assign LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_mx0w0 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      dma_read_chnl_rsci_idat_mxwt, LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_1);
  assign LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0 = MUX_v_32_2_2(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d_mxwt,
      LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1, LOAD_LOOP_for_if_2_for_for_asn_126_itm_2);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_61_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_29_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_0_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_0_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_60_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_28_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_1_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_1_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_59_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_27_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_2_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_2_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_58_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_26_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_3_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_3_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_57_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_25_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_4_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_4_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_56_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_24_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_5_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_5_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_55_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_23_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_6_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_6_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_54_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_22_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_7_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_7_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_53_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_21_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_8_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_8_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_52_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_20_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_9_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_9_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_51_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_19_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_10_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_10_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_50_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_18_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_11_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_11_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_49_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_17_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_12_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_12_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_48_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_16_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_13_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_13_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_47_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_15_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_14_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_14_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_46_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_14_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_15_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_15_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_45_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_13_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_16_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_16_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_44_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_12_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_17_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_17_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_43_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_11_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_18_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_18_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_42_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_10_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_19_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_19_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_41_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_9_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_20_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_20_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_40_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_8_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_21_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_21_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_39_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_7_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_22_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_22_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_38_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_6_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_23_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_23_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_37_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_5_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_24_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_24_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_36_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_4_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_25_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_25_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_35_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_3_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_26_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_26_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_34_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_2_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_27_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_27_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_33_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_1_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_28_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_28_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_32_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_0_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_29_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_29_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_31_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_31_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_5_30_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_4_30_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_31_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_15_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_30_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_14_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_0_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_0_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_1_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_1_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_2_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_2_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_3_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_3_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_4_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_4_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_5_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_5_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_6_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_6_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_7_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_7_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_8_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_8_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_9_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_9_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_10_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_10_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_11_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_11_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_12_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_12_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_13_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_13_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_14_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_14_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_15_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_15_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_16_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_0_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_17_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_1_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_18_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_2_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_19_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_3_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_20_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_4_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_21_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_5_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_22_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_6_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_23_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_7_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_24_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_8_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_25_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_9_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_26_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_10_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_27_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_11_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_28_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_12_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_4_29_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_3_13_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_14_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_6_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_15_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_7_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_0_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_0_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_1_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_1_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_2_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_2_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_3_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_3_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_4_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_4_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_5_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_5_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_6_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_6_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_7_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_7_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_8_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_0_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_9_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_1_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_10_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_2_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_11_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_3_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_12_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_4_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_3_13_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_2_5_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_6_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_7_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_0_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_1_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_2_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_3_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]));
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_4_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign LOAD_LOOP_for_if_2_for_for_and_stg_2_5_sva_1 = LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1 = MUX_v_5_2_2(5'b00000, LOAD_LOOP_for_k_5_0_lpi_2_4_0,
      lfst_exit_LOAD_LOOP_sva);
  assign nl_operator_8_false_1_acc_tmp = conv_u2s_8_9(conf_info_crt_sva_231_0[103:96])
      + 9'b111111111;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[8:0];
  assign LOAD_LOOP_for_if_for_for_if_nor_cse_sva_1 = ~((operator_8_false_1_acc_tmp[7:3]!=5'b00000));
  assign nl_operator_8_false_4_acc_nl = ({1'b1 , LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1})
      + 4'b0001;
  assign operator_8_false_4_acc_nl = nl_operator_8_false_4_acc_nl[3:0];
  assign operator_8_false_4_acc_itm_3_1 = readslicef_4_1_3(operator_8_false_4_acc_nl);
  assign nl_LOAD_BATCH_LOOP_acc_tmp = conv_u2u_4_5(LOAD_BATCH_LOOP_b_4_0_sva_3_0)
      + 5'b00001;
  assign LOAD_BATCH_LOOP_acc_tmp = nl_LOAD_BATCH_LOOP_acc_tmp[4:0];
  assign LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_nor_tmp = ~((~((LOAD_BATCH_LOOP_b_4_0_sva_3_0
      == (operator_8_false_8_acc_psp_sva_1[3:0])) & (operator_8_false_8_acc_psp_sva_1[7:4]==4'b0000)))
      | (operator_8_false_8_acc_psp_sva_1[8]));
  assign nl_operator_8_false_8_acc_psp_sva_1 = conv_u2s_8_9(conf_info_crt_sva_231_0[231:224])
      + 9'b111111111;
  assign operator_8_false_8_acc_psp_sva_1 = nl_operator_8_false_8_acc_psp_sva_1[8:0];
  assign nl_LOAD_LOOP_acc_tmp = conv_u2u_5_6(LOAD_LOOP_fl_5_0_sva_4_0) + 6'b000001;
  assign LOAD_LOOP_acc_tmp = nl_LOAD_LOOP_acc_tmp[5:0];
  assign LOAD_LOOP_if_equal_tmp = LOAD_LOOP_fl_5_0_sva_4_0 == (operator_8_false_7_acc_tmp[4:0]);
  assign exit_LOAD_LOOP_sva_3 = ~((~(LOAD_LOOP_if_equal_tmp & (operator_8_false_7_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_7_acc_tmp[8]));
  assign nl_operator_8_false_7_acc_tmp = conv_u2s_8_9(conf_info_crt_sva_231_0[71:64])
      + 9'b111111111;
  assign operator_8_false_7_acc_tmp = nl_operator_8_false_7_acc_tmp[8:0];
  assign nl_LOAD_LOOP_for_acc_2_tmp = conv_u2u_5_6(LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1)
      + 6'b000001;
  assign LOAD_LOOP_for_acc_2_tmp = nl_LOAD_LOOP_for_acc_2_tmp[5:0];
  assign LOAD_LOOP_for_if_3_equal_tmp = LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1 == (operator_8_false_6_acc_tmp[4:0]);
  assign LOAD_LOOP_for_if_2_for_mux_5_nl = MUX_s_1_2_2(or_810_cse, exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm,
      and_dcpl_778);
  assign exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_3 = LOAD_LOOP_for_if_2_for_mux_5_nl
      & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0;
  assign nl_LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_1_nl = conv_u2u_8_9({(~ n_w_in_acc_psp_sva)
      , (~ (conf_info_crt_sva_231_0[192]))}) + conv_u2u_8_9(pad_sva) + 9'b000000001;
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_1_nl = nl_LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_1_nl[8:0];
  assign nl_LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_nl = conv_u2u_9_10(LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_1_nl)
      + conv_s2u_9_10({4'b1000 , LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1});
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_nl = nl_LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_nl[9:0];
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_itm_9_1 = readslicef_10_1_9(LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_nl);
  assign nl_LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_1_nl = conv_u2u_8_9({(~ n_h_in_acc_psp_sva)
      , (~ (conf_info_crt_sva_231_0[160]))}) + conv_u2u_8_9(pad_sva) + 9'b000000001;
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_1_nl = nl_LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_1_nl[8:0];
  assign nl_LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_nl = conv_u2u_9_10(LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_1_nl)
      + conv_s2u_9_10({4'b1000 , LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1});
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_nl = nl_LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_nl[9:0];
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_itm_9_1 = readslicef_10_1_9(LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_nl);
  assign nl_operator_8_false_6_acc_tmp = conv_u2s_8_9(conf_info_crt_sva_231_0[135:128])
      + 9'b111111111;
  assign operator_8_false_6_acc_tmp = nl_operator_8_false_6_acc_tmp[8:0];
  assign nl_operator_8_false_5_acc_nl = conv_u2s_4_5(LOAD_LOOP_for_if_2_for_row_4_0_sva_1_mx0w1[4:1])
      + 5'b10111;
  assign operator_8_false_5_acc_nl = nl_operator_8_false_5_acc_nl[4:0];
  assign operator_8_false_5_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_5_acc_nl);
  assign nl_operator_8_false_5_acc_psp_sva_1 = conv_u2s_8_9({n_w_in_acc_psp_sva ,
      (conf_info_crt_sva_231_0[192])}) + 9'b111111111;
  assign operator_8_false_5_acc_psp_sva_1 = nl_operator_8_false_5_acc_psp_sva_1[8:0];
  assign nl_operator_8_false_4_acc_psp_sva_1 = conv_u2s_8_9({n_h_in_acc_psp_sva ,
      (conf_info_crt_sva_231_0[160])}) + 9'b111111111;
  assign operator_8_false_4_acc_psp_sva_1 = nl_operator_8_false_4_acc_psp_sva_1[8:0];
  assign LOAD_LOOP_for_if_for_for_and_stg_4_16_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_0_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]);
  assign LOAD_LOOP_for_if_for_for_and_stg_4_0_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_0_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_15_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_15_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_1_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_1_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_14_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_14_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_2_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_2_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_13_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_13_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_3_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_3_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_12_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_12_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_4_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_4_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_11_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_11_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_5_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_5_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_10_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_10_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_6_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_6_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_9_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_9_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_7_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_7_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_4_8_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_3_8_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_15_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_7_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_1_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_1_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_14_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_6_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_2_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_2_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_13_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_5_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_3_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_3_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_12_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_4_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_4_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_4_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_11_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_3_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_5_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_5_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_10_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_2_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_6_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_6_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_9_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_1_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_7_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_7_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_3_8_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_0_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign LOAD_LOOP_for_if_for_for_and_stg_3_0_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_2_0_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign LOAD_LOOP_for_if_for_for_and_stg_2_1_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_1_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign LOAD_LOOP_for_if_for_for_and_stg_2_2_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_2_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign LOAD_LOOP_for_if_for_for_and_stg_2_3_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_3_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign LOAD_LOOP_for_if_for_for_and_stg_2_4_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_0_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign LOAD_LOOP_for_if_for_for_and_stg_2_5_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_1_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign LOAD_LOOP_for_if_for_for_and_stg_2_6_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_2_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign LOAD_LOOP_for_if_for_for_and_stg_2_7_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_3_sva_1
      & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign LOAD_LOOP_for_if_for_for_and_stg_2_0_sva_1 = LOAD_LOOP_for_if_for_for_and_stg_1_0_sva_1
      & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign LOAD_LOOP_for_if_for_for_and_stg_1_1_sva_1 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]==2'b01);
  assign LOAD_LOOP_for_if_for_for_and_stg_1_2_sva_1 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]==2'b10);
  assign LOAD_LOOP_for_if_for_for_and_stg_1_3_sva_1 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]==2'b11);
  assign LOAD_LOOP_for_if_for_for_and_stg_1_0_sva_1 = ~((LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]!=2'b00));
  assign exitL_exit_LOAD_CTRL_LOOP2_lpi_2_dfm_1 = dma_read_ctrl_rsci_irdy_mxwt |
      (~ LOAD_LOOP_for_asn_6_itm_1);
  assign LOAD_LOOP_for_if_2_for_and_181_cse_1 = exitL_exit_LOAD_CTRL_LOOP2_lpi_2_dfm_1
      & LOAD_LOOP_for_if_2_for_equal_tmp_1_1;
  assign LOAD_LOOP_for_if_2_for_and_180_cse_1 = (~ exitL_exit_LOAD_CTRL_LOOP2_lpi_2_dfm_1)
      & LOAD_LOOP_for_if_2_for_equal_tmp_1_1;
  assign LOAD_LOOP_for_if_2_for_and_178_m1c_1 = (~ exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_1)
      & LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
  assign LOAD_LOOP_for_if_2_for_for_and_251_tmp_1 = (~ exit_LOAD_LOOP_for_if_2_for_sva_1_1)
      & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_1;
  assign LOAD_LOOP_for_if_2_for_and_176_m1c_1 = (~ exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_1)
      & LOAD_LOOP_for_if_2_for_equal_tmp_1;
  assign LOAD_LOOP_for_if_for_for_and_tmp_1 = (~ exit_LOAD_LOOP_for_if_for_sva_1_1)
      & exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_1;
  assign LOAD_LOOP_for_if_2_for_for_and_250_tmp_1 = LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_1
      & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_1;
  assign LOAD_LOOP_for_if_2_for_and_195_ssc_1 = exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_1
      & LOAD_LOOP_for_if_2_for_equal_tmp_1;
  assign LOAD_LOOP_mux_1_nl = MUX_s_1_2_2(exit_LOAD_LOOP_lpi_2_dfm_1_mx0w0, exit_LOAD_LOOP_lpi_2_dfm_1,
      or_dcpl_150);
  assign exit_LOAD_LOOP_lpi_2_dfm_4 = LOAD_LOOP_mux_1_nl & exit_LOAD_LOOP_for_lpi_2_dfm_3_mx0w0;
  assign LOAD_LOOP_for_LOAD_LOOP_nand_cse = ~(lfst_exit_LOAD_LOOP_for_1_lpi_2 & lfst_exit_LOAD_LOOP_sva);
  assign LOAD_LOOP_for_if_2_for_mux_22_nl = MUX_s_1_2_2(exitL_exit_LOAD_LOOP_for_if_2_for_sva_1_mx0w0,
      exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2, or_75_cse);
  assign exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1 = LOAD_LOOP_for_if_2_for_mux_22_nl
      | LOAD_LOOP_for_LOAD_LOOP_nand_cse;
  assign LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1 = buf_linear_rsci_bawt | (~(LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3
      & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3 & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2
      & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0==2'b00) & LOAD_BATCH_LOOP_stage_v_3));
  assign operator_8_false_operator_8_false_nor_cse_sva_1 = ~((LOAD_LOOP_fl_5_0_sva_4_0!=5'b00000));
  assign LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_and_cse_1 = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1[0])
      & (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1[1])));
  assign LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_nor_1_cse_1 = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1
      | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1!=2'b00));
  assign nl_operator_8_false_1_acc_4_nl = conv_u2u_1_2(~ (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[1]))
      + conv_u2u_1_2(LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[2]) + conv_u2u_1_2(~
      (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[3]));
  assign operator_8_false_1_acc_4_nl = nl_operator_8_false_1_acc_4_nl[1:0];
  assign nl_operator_8_false_1_acc_psp_sva_1 = conv_u2s_2_3(operator_8_false_1_acc_4_nl)
      + conv_s2s_2_3({1'b1 , (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[0])}) + conv_u2s_1_3(LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[4]);
  assign operator_8_false_1_acc_psp_sva_1 = nl_operator_8_false_1_acc_psp_sva_1[2:0];
  assign nl_operator_8_false_3_acc_2_nl = ({(~ (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[2]))
      , 2'b00}) + conv_u2u_2_3(LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[4:3]) + conv_u2u_1_3(LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[2]);
  assign operator_8_false_3_acc_2_nl = nl_operator_8_false_3_acc_2_nl[2:0];
  assign nl_operator_8_false_3_acc_psp_sva_1 = conv_u2s_3_4(operator_8_false_3_acc_2_nl)
      + conv_s2s_3_4({1'b1 , (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[1:0])});
  assign operator_8_false_3_acc_psp_sva_1 = nl_operator_8_false_3_acc_psp_sva_1[3:0];
  assign nl_LOAD_LOOP_for_if_2_for_for_acc_2_psp_1 = (LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1[4:1])
      + conv_u2u_3_4(LOAD_LOOP_for_if_2_for_for_row_norm_2_0_lpi_2_dfm_1);
  assign LOAD_LOOP_for_if_2_for_for_acc_2_psp_1 = nl_LOAD_LOOP_for_if_2_for_for_acc_2_psp_1[3:0];
  assign nl_operator_8_false_1_acc_3_nl = conv_u2u_1_2(z_out_7[0]) + conv_u2u_1_2(z_out_7[1]);
  assign operator_8_false_1_acc_3_nl = nl_operator_8_false_1_acc_3_nl[1:0];
  assign nl_operator_8_false_3_operator_8_false_3_acc_nl = conv_s2u_1_3(z_out_9[2])
      + z_out_9;
  assign operator_8_false_3_operator_8_false_3_acc_nl = nl_operator_8_false_3_operator_8_false_3_acc_nl[2:0];
  assign LOAD_LOOP_for_if_2_for_for_switch_lp_LOAD_LOOP_for_if_2_for_for_switch_lp_and_3_nl
      = (conf_info_crt_sva_231_0[103:96]==8'b00000111);
  assign LOAD_LOOP_for_if_2_for_for_switch_lp_mux1h_4_nl = MUX1HOT_v_3_3_2(({1'b0
      , operator_8_false_1_acc_3_nl}), z_out_7, operator_8_false_3_operator_8_false_3_acc_nl,
      {(~ (conf_info_crt_sva_231_0[98])) , (~ (conf_info_crt_sva_231_0[97])) , LOAD_LOOP_for_if_2_for_for_switch_lp_LOAD_LOOP_for_if_2_for_for_switch_lp_and_3_nl});
  assign LOAD_LOOP_for_if_2_for_for_switch_lp_nand_nl = ~((conf_info_crt_sva_231_0[103:96]==8'b00000001));
  assign LOAD_LOOP_for_if_2_for_for_row_norm_2_0_lpi_2_dfm_1 = MUX_v_3_2_2(3'b000,
      LOAD_LOOP_for_if_2_for_for_switch_lp_mux1h_4_nl, LOAD_LOOP_for_if_2_for_for_switch_lp_nand_nl);
  assign LOAD_BATCH_LOOP_and_4_tmp = LOAD_BATCH_LOOP_stage_v & (~(LOAD_BATCH_LOOP_stage_v_1
      & (~ LOAD_BATCH_LOOP_and_3_tmp))) & LOAD_BATCH_LOOP_stage_0_1 & (plm_kernel_rsci_bawt
      | (~(exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2 & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1])
      & (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0])))
      & LOAD_BATCH_LOOP_stage_v_2))) & (LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt
      | (~(LOAD_LOOP_for_if_2_for_for_asn_itm_2 & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2
      & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0==2'b00) & LOAD_BATCH_LOOP_stage_v_2)))
      & LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1;
  assign LOAD_BATCH_LOOP_and_3_tmp = LOAD_BATCH_LOOP_stage_v_1 & (~(LOAD_BATCH_LOOP_stage_v_2
      & or_dcpl_135)) & LOAD_BATCH_LOOP_stage_0_2 & (dma_read_ctrl_rsci_bawt | (~(((lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0])
      & (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]))))
      | (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0!=2'b00))))))
      & (dma_read_chnl_rsci_bawt | (~((lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1])
      & (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]))))))
      & (dma_read_ctrl_rsci_bawt | (~(LOAD_LOOP_for_asn_2_itm_1 & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0==2'b11)
      & (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2)))) & (dma_read_chnl_rsci_bawt
      | (~(LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st_1 & LOAD_LOOP_for_if_2_for_for_asn_itm_1
      & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0==2'b00))))
      & LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1;
  assign or_tmp_4 = (~ LOAD_BATCH_LOOP_stage_v_3) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0!=2'b00)
      | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2) | (~ exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3)
      | (~ LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3) | buf_linear_rsci_bawt;
  assign or_9_cse = (~ LOAD_LOOP_for_if_2_for_for_asn_itm_2) | LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt;
  assign or_41_cse = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0!=2'b00);
  assign or_42_cse = (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]))
      | plm_kernel_rsci_bawt | (~ exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign or_44_cse = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2) | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00);
  assign and_3266_cse = lfst_exit_LOAD_LOOP_sva & lfst_exit_LOAD_LOOP_for_1_lpi_2;
  assign or_tmp_57 = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2 | (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]))
      | plm_kernel_rsci_bawt | (~ exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign and_tmp_12 = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 & (~(LOAD_LOOP_for_asn_6_itm_1
      & (~ dma_read_ctrl_rsci_irdy_mxwt)));
  assign or_tmp_90 = LOAD_BATCH_LOOP_stage_0 | (~ or_654_cse);
  assign mux_1110_nl = MUX_s_1_2_2(or_tmp_90, (~ or_654_cse), exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign mux_1109_nl = MUX_s_1_2_2(or_tmp_90, mux_1110_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_tmp_52 = MUX_s_1_2_2(mux_1109_nl, or_tmp_90, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign nor_37_cse = ~(LOAD_BATCH_LOOP_asn_itm_1 | (~ LOAD_BATCH_LOOP_and_3_tmp));
  assign or_93_cse = (~ LOAD_LOOP_for_if_2_for_equal_tmp_2_1) | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2)
      | LOAD_LOOP_for_if_2_for_or_tmp_1;
  assign or_101_cse = (~((~ LOAD_LOOP_for_if_2_for_equal_tmp_2_1) | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2))
      | LOAD_LOOP_for_if_2_for_or_tmp_1;
  assign nor_tmp_50 = ~(dma_read_ctrl_rsci_irdy_mxwt | (~ LOAD_LOOP_for_asn_6_itm_1));
  assign mux_74_nl = MUX_s_1_2_2(or_tmp_90, (~ or_654_cse), exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign mux_75_nl = MUX_s_1_2_2(or_tmp_90, mux_74_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_1101_nl = MUX_s_1_2_2(mux_75_nl, or_tmp_90, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign mux_79_nl = MUX_s_1_2_2(or_tmp_90, mux_1101_nl, and_3192_cse);
  assign mux_1140_nl = MUX_s_1_2_2(or_tmp_90, (~ or_654_cse), exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign mux_1139_nl = MUX_s_1_2_2(or_tmp_90, mux_1140_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_1100_nl = MUX_s_1_2_2(mux_1139_nl, or_tmp_90, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign mux_78_nl = MUX_s_1_2_2(or_tmp_90, mux_1100_nl, nor_225_cse);
  assign mux_80_nl = MUX_s_1_2_2(mux_79_nl, mux_78_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_51_nl = MUX_s_1_2_2(or_tmp_90, (~ or_654_cse), exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign mux_52_nl = MUX_s_1_2_2(or_tmp_90, mux_51_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_1108_nl = MUX_s_1_2_2(mux_52_nl, or_tmp_90, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign mux_54_nl = MUX_s_1_2_2(or_tmp_90, mux_1108_nl, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_tmp_80 = MUX_s_1_2_2(mux_80_nl, mux_54_nl, or_750_cse);
  assign mux_1120_nl = MUX_s_1_2_2(or_tmp_90, (~ or_654_cse), exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign mux_1119_nl = MUX_s_1_2_2(or_tmp_90, mux_1120_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_316_nl = MUX_s_1_2_2(mux_1119_nl, or_tmp_90, or_755_cse);
  assign mux_83_nl = MUX_s_1_2_2(mux_tmp_52, mux_tmp_80, or_101_cse);
  assign mux_82_nl = MUX_s_1_2_2(mux_tmp_52, mux_tmp_80, or_93_cse);
  assign mux_84_nl = MUX_s_1_2_2(mux_83_nl, mux_82_nl, or_44_cse);
  assign mux_86_nl = MUX_s_1_2_2(mux_316_nl, mux_84_nl, nor_37_cse);
  assign and_3236_nl = or_2860_cse & lfst_exit_LOAD_LOOP_for_1_lpi_2 & lfst_exit_LOAD_LOOP_sva
      & LOAD_BATCH_LOOP_and_4_tmp;
  assign mux_87_nl = MUX_s_1_2_2(or_tmp_90, mux_86_nl, and_3236_nl);
  assign mux_88_nl = MUX_s_1_2_2(or_tmp_90, mux_87_nl, or_513_cse);
  assign mux_89_nl = MUX_s_1_2_2(or_tmp_90, mux_88_nl, or_810_cse);
  assign and_dcpl_24 = (~ mux_89_nl) & (~(LOAD_BATCH_LOOP_stage_0_2 | LOAD_BATCH_LOOP_stage_0_3))
      & LOAD_BATCH_LOOP_stage_v_3 & (~ LOAD_BATCH_LOOP_stage_0_1);
  assign nor_tmp_54 = dma_read_ctrl_rsci_irdy_mxwt & LOAD_LOOP_for_if_2_for_equal_tmp_1_1;
  assign or_tmp_148 = (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1])))
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign and_tmp_17 = or_75_cse & or_tmp_148;
  assign or_tmp_151 = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign nor_55_cse = ~(LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (~ (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1])));
  assign or_180_nl = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1])
      | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign mux_90_nl = MUX_s_1_2_2(or_180_nl, or_tmp_151, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_177_nl = nor_55_cse | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign mux_91_nl = MUX_s_1_2_2(mux_90_nl, or_177_nl, LOAD_LOOP_for_if_2_for_or_tmp_1);
  assign mux_tmp_91 = MUX_s_1_2_2((~ mux_91_nl), or_tmp_148, or_75_cse);
  assign mux_tmp_93 = MUX_s_1_2_2(mux_tmp_91, and_tmp_17, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign and_dcpl_28 = and_3266_cse & LOAD_BATCH_LOOP_and_4_tmp & LOAD_LOOP_for_asn_sft_lpi_2;
  assign or_tmp_154 = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2) | LOAD_LOOP_for_if_2_for_or_tmp_1;
  assign mux_tmp_103 = MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_mux_11_itm_1, mux_335_cse,
      LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign or_192_nl = (~((~((lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b10)))
      | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2)) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign mux_107_cse = MUX_s_1_2_2(or_tmp_148, or_192_nl, LOAD_LOOP_for_asn_sft_lpi_2);
  assign nor_tmp_63 = ~(LOAD_LOOP_for_if_2_for_or_tmp_1 | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2));
  assign mux_1148_nl = MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_equal_tmp_1_1, nor_tmp_54,
      LOAD_LOOP_for_asn_2_itm_1);
  assign mux_1147_nl = MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_equal_tmp_1_1, mux_1148_nl,
      LOAD_LOOP_for_asn_6_itm_1);
  assign mux_tmp_109 = MUX_s_1_2_2(mux_1147_nl, LOAD_LOOP_for_if_2_for_equal_tmp_1_1,
      or_750_cse);
  assign nand_24_cse = ~(LOAD_LOOP_for_if_2_for_and_195_ssc_1 & (~ mux_tmp_109));
  assign nor_tmp_67 = ~(LOAD_LOOP_for_if_2_for_or_tmp_1 | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2));
  assign or_197_cse = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | mux_tmp_109;
  assign and_dcpl_33 = ~((LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[0]) | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign and_dcpl_34 = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]) &
      (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2);
  assign and_dcpl_35 = and_dcpl_34 & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1]));
  assign and_dcpl_36 = and_dcpl_35 & and_dcpl_33;
  assign and_dcpl_38 = ~((LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]!=2'b00)
      | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]));
  assign and_dcpl_39 = LOAD_BATCH_LOOP_and_3_tmp & exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_1;
  assign and_dcpl_40 = and_dcpl_39 & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]));
  assign and_dcpl_41 = and_dcpl_40 & and_dcpl_38;
  assign and_dcpl_44 = and_dcpl_39 & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]))
      & and_dcpl_34;
  assign or_dcpl_29 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]!=2'b00);
  assign or_dcpl_30 = or_dcpl_29 | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign or_dcpl_31 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4:3]!=2'b00);
  assign or_dcpl_32 = or_dcpl_31 | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
  assign or_dcpl_34 = (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]))
      | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2;
  assign and_dcpl_46 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[0]) & (~
      (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign and_dcpl_47 = and_dcpl_35 & and_dcpl_46;
  assign or_dcpl_38 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]!=2'b01);
  assign or_dcpl_39 = or_dcpl_38 | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign and_dcpl_50 = and_dcpl_34 & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1]);
  assign and_dcpl_51 = and_dcpl_50 & and_dcpl_33;
  assign or_dcpl_41 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]!=2'b10);
  assign or_dcpl_42 = or_dcpl_41 | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign and_dcpl_54 = and_dcpl_50 & and_dcpl_46;
  assign or_dcpl_44 = ~((LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[1:0]==2'b11));
  assign or_dcpl_45 = or_dcpl_44 | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign and_dcpl_57 = (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[0])) &
      (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign and_dcpl_58 = and_dcpl_35 & and_dcpl_57;
  assign or_dcpl_47 = or_dcpl_29 | (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign and_dcpl_61 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[0]) & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]);
  assign and_dcpl_62 = and_dcpl_35 & and_dcpl_61;
  assign or_dcpl_49 = or_dcpl_38 | (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign and_dcpl_65 = and_dcpl_50 & and_dcpl_57;
  assign or_dcpl_51 = or_dcpl_41 | (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign and_dcpl_68 = and_dcpl_50 & and_dcpl_61;
  assign or_dcpl_53 = or_dcpl_44 | (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[2]));
  assign and_dcpl_71 = and_dcpl_39 & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[3]);
  assign and_dcpl_72 = and_dcpl_71 & and_dcpl_38;
  assign or_dcpl_55 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4:3]!=2'b01);
  assign or_dcpl_56 = or_dcpl_55 | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
  assign and_dcpl_90 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01)
      & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]));
  assign and_dcpl_91 = and_dcpl_40 & and_dcpl_90;
  assign or_dcpl_65 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[4:3]!=2'b10);
  assign or_dcpl_66 = or_dcpl_65 | (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
  assign and_dcpl_108 = and_dcpl_71 & and_dcpl_90;
  assign or_dcpl_76 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:3]!=3'b011);
  assign and_dcpl_126 = (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b10)
      & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]));
  assign and_dcpl_127 = and_dcpl_40 & and_dcpl_126;
  assign or_dcpl_85 = or_dcpl_31 | (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
  assign and_dcpl_144 = and_dcpl_71 & and_dcpl_126;
  assign or_dcpl_94 = or_dcpl_55 | (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
  assign or_dcpl_103 = or_dcpl_65 | (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
  assign and_dcpl_166 = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00));
  assign and_dcpl_167 = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b00));
  assign and_dcpl_168 = and_dcpl_167 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign and_dcpl_169 = and_dcpl_168 & and_dcpl_166;
  assign and_dcpl_170 = LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_2
      & LOAD_BATCH_LOOP_stage_0_3;
  assign and_dcpl_172 = (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]))
      & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2;
  assign and_dcpl_173 = and_dcpl_172 & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_2;
  assign and_dcpl_174 = and_dcpl_173 & and_dcpl_170 & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1;
  assign and_dcpl_176 = LOAD_BATCH_LOOP_stage_v_2 & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]));
  assign and_dcpl_178 = or_tmp_4 & and_dcpl_176 & or_9_cse;
  assign and_dcpl_182 = and_dcpl_176 & and_dcpl_172;
  assign and_dcpl_183 = and_dcpl_182 & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_2
      & LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_2 & LOAD_BATCH_LOOP_stage_0_3;
  assign not_tmp_118 = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 | (~ or_tmp_4));
  assign and_dcpl_186 = (~ LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_bawt) & LOAD_LOOP_for_if_2_for_for_asn_itm_2;
  assign and_dcpl_188 = and_dcpl_173 & and_dcpl_170 & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1;
  assign not_tmp_124 = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 | (~ or_tmp_4));
  assign and_dcpl_194 = and_dcpl_173 & and_dcpl_170 & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1;
  assign not_tmp_125 = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 | (~ or_tmp_4));
  assign and_dcpl_200 = and_dcpl_173 & and_dcpl_170 & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1;
  assign not_tmp_126 = ~(LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 | (~ or_tmp_4));
  assign and_dcpl_205 = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b01);
  assign and_dcpl_206 = and_dcpl_168 & and_dcpl_205;
  assign and_dcpl_223 = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b10);
  assign and_dcpl_224 = and_dcpl_168 & and_dcpl_223;
  assign and_dcpl_241 = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11);
  assign and_dcpl_242 = and_dcpl_168 & and_dcpl_241;
  assign and_dcpl_259 = and_dcpl_167 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign and_dcpl_260 = and_dcpl_259 & and_dcpl_166;
  assign and_dcpl_277 = and_dcpl_259 & and_dcpl_205;
  assign and_dcpl_294 = and_dcpl_259 & and_dcpl_223;
  assign and_dcpl_311 = and_dcpl_259 & and_dcpl_241;
  assign and_dcpl_328 = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b01);
  assign and_dcpl_329 = and_dcpl_328 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign and_dcpl_330 = and_dcpl_329 & and_dcpl_166;
  assign and_dcpl_347 = and_dcpl_329 & and_dcpl_205;
  assign and_dcpl_364 = and_dcpl_329 & and_dcpl_223;
  assign and_dcpl_381 = and_dcpl_329 & and_dcpl_241;
  assign and_dcpl_398 = and_dcpl_328 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign and_dcpl_399 = and_dcpl_398 & and_dcpl_166;
  assign and_dcpl_416 = and_dcpl_398 & and_dcpl_205;
  assign and_dcpl_433 = and_dcpl_398 & and_dcpl_223;
  assign and_dcpl_450 = and_dcpl_398 & and_dcpl_241;
  assign and_dcpl_467 = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b10);
  assign and_dcpl_468 = and_dcpl_467 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign and_dcpl_469 = and_dcpl_468 & and_dcpl_166;
  assign not_tmp_127 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1)) & or_tmp_4;
  assign not_tmp_128 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1)) & or_tmp_4;
  assign not_tmp_129 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1)) & or_tmp_4;
  assign not_tmp_130 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1)) & or_tmp_4;
  assign and_dcpl_486 = and_dcpl_468 & and_dcpl_205;
  assign and_dcpl_503 = and_dcpl_468 & and_dcpl_223;
  assign and_dcpl_520 = and_dcpl_468 & and_dcpl_241;
  assign and_dcpl_537 = and_dcpl_467 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign and_dcpl_538 = and_dcpl_537 & and_dcpl_166;
  assign and_dcpl_555 = and_dcpl_537 & and_dcpl_205;
  assign and_dcpl_572 = and_dcpl_537 & and_dcpl_223;
  assign and_dcpl_589 = and_dcpl_537 & and_dcpl_241;
  assign and_dcpl_606 = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b11);
  assign and_dcpl_607 = and_dcpl_606 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]));
  assign and_dcpl_608 = and_dcpl_607 & and_dcpl_166;
  assign not_tmp_131 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1)) & or_tmp_4;
  assign not_tmp_132 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1)) & or_tmp_4;
  assign not_tmp_133 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1)) & or_tmp_4;
  assign not_tmp_134 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1)) & or_tmp_4;
  assign and_dcpl_625 = and_dcpl_607 & and_dcpl_205;
  assign and_dcpl_642 = and_dcpl_607 & and_dcpl_223;
  assign and_dcpl_659 = and_dcpl_607 & and_dcpl_241;
  assign and_dcpl_676 = and_dcpl_606 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign and_dcpl_677 = and_dcpl_676 & and_dcpl_166;
  assign not_tmp_135 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1)) & or_tmp_4;
  assign not_tmp_136 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1)) & or_tmp_4;
  assign not_tmp_137 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1)) & or_tmp_4;
  assign not_tmp_138 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1)) & or_tmp_4;
  assign and_dcpl_694 = and_dcpl_676 & and_dcpl_205;
  assign and_dcpl_711 = and_dcpl_676 & and_dcpl_223;
  assign and_dcpl_728 = and_dcpl_676 & and_dcpl_241;
  assign and_dcpl_738 = LOAD_BATCH_LOOP_and_3_tmp & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]));
  assign and_dcpl_739 = and_dcpl_738 & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]));
  assign and_dcpl_752 = and_3266_cse & LOAD_BATCH_LOOP_and_4_tmp;
  assign or_tmp_325 = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | (~ and_tmp_12);
  assign nor_tmp_101 = lfst_exit_LOAD_LOOP_for_1_lpi_2 & lfst_exit_LOAD_LOOP_sva
      & LOAD_BATCH_LOOP_and_4_tmp;
  assign mux_260_nl = MUX_s_1_2_2((~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2),
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]);
  assign mux_tmp_260 = MUX_s_1_2_2(or_dcpl_34, mux_260_nl, and_3198_cse);
  assign nand_tmp_29 = ~(LOAD_LOOP_for_if_2_for_and_195_ssc_1 & (~ mux_tmp_260));
  assign or_tmp_340 = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]) |
      mux_tmp_260;
  assign and_3239_nl = dma_read_ctrl_rsci_irdy_mxwt & LOAD_LOOP_for_asn_2_itm_1 &
      (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]) & (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2);
  assign mux_278_nl = MUX_s_1_2_2((~ or_dcpl_34), and_3239_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign and_tmp_22 = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 & mux_278_nl;
  assign nor_113_cse = ~(nor_tmp_67 | (~ (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1])));
  assign or_461_itm = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | LOAD_LOOP_for_if_2_for_equal_tmp_2_1
      | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0]);
  assign mux_1156_nl = MUX_s_1_2_2(mux_1159_itm, or_tmp_340, or_461_itm);
  assign mux_282_nl = MUX_s_1_2_2(mux_1156_nl, or_tmp_340, LOAD_BATCH_LOOP_asn_itm_1);
  assign nand_tmp_32 = ~(LOAD_BATCH_LOOP_and_3_tmp & (~ mux_282_nl));
  assign or_468_nl = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 | (~ mux_tmp_260);
  assign mux_tmp_284 = MUX_s_1_2_2(or_468_nl, and_tmp_22, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]);
  assign or_470_nl = (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1]) | mux_tmp_284;
  assign nand_33_nl = ~((LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1]) & (~ mux_tmp_284));
  assign mux_286_nl = MUX_s_1_2_2(or_470_nl, nand_33_nl, nor_tmp_67);
  assign mux_287_nl = MUX_s_1_2_2(mux_286_nl, mux_tmp_284, LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0]);
  assign or_469_nl = nor_tmp_63 | mux_tmp_284;
  assign mux_288_nl = MUX_s_1_2_2(mux_287_nl, or_469_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_1157_itm = MUX_s_1_2_2((~ mux_288_nl), or_tmp_340, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign mux_290_nl = MUX_s_1_2_2(mux_1157_itm, or_tmp_340, LOAD_BATCH_LOOP_asn_itm_1);
  assign nand_tmp_34 = ~(LOAD_BATCH_LOOP_and_3_tmp & (~ mux_290_nl));
  assign or_tmp_352 = or_75_cse | (~ mux_1157_itm);
  assign and_dcpl_764 = and_dcpl_176 & exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2
      & plm_kernel_rsci_bawt & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1])
      & (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2) & LOAD_BATCH_LOOP_stage_0_3;
  assign and_dcpl_772 = (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0[0]))
      & lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2 & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0[1]))
      & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3 & LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3
      & buf_linear_rsci_bawt & LOAD_BATCH_LOOP_stage_v_3;
  assign or_dcpl_122 = (~ LOAD_BATCH_LOOP_stage_v_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign or_dcpl_128 = (~ LOAD_BATCH_LOOP_and_3_tmp) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]);
  assign or_dcpl_129 = or_dcpl_128 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[1]);
  assign or_tmp_388 = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2) | LOAD_LOOP_for_if_2_for_or_tmp_1;
  assign mux_17_nl = MUX_s_1_2_2(or_42_cse, or_41_cse, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign mux_332_nl = MUX_s_1_2_2(mux_17_nl, or_tmp_57, or_9_cse);
  assign and_tmp_25 = or_tmp_4 & mux_332_nl;
  assign or_dcpl_135 = ~(and_tmp_25 & LOAD_BATCH_LOOP_stage_v_2 & LOAD_BATCH_LOOP_stage_0_3);
  assign or_dcpl_136 = LOAD_LOOP_for_LOAD_LOOP_nand_cse | (~ LOAD_BATCH_LOOP_and_4_tmp);
  assign and_dcpl_778 = (~ LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_if_1_LOAD_LOOP_for_if_2_for_for_if_1_nor_tmp)
      & operator_8_false_6_acc_itm_4_1;
  assign or_dcpl_146 = ~((~ and_dcpl_778) & lfst_exit_LOAD_LOOP_for_1_lpi_2 & lfst_exit_LOAD_LOOP_sva
      & LOAD_BATCH_LOOP_and_4_tmp);
  assign and_dcpl_779 = operator_8_false_5_acc_itm_4_1 & (~ LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_1_LOAD_LOOP_for_if_2_for_if_1_nor_tmp);
  assign or_tmp_408 = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | (~ or_2860_cse);
  assign or_tmp_409 = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | (~ or_2860_cse);
  assign mux_tmp_336 = MUX_s_1_2_2(or_tmp_409, or_tmp_408, or_75_cse);
  assign or_559_nl = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2) | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00)
      | or_tmp_409;
  assign nand_36_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 & (~ or_tmp_409));
  assign mux_338_nl = MUX_s_1_2_2(or_559_nl, nand_36_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_560_nl = LOAD_LOOP_for_if_2_for_or_tmp_1 | mux_338_nl;
  assign mux_tmp_338 = MUX_s_1_2_2(or_560_nl, or_tmp_408, or_75_cse);
  assign mux_tmp_340 = MUX_s_1_2_2(mux_tmp_338, mux_tmp_336, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_340_nl = MUX_s_1_2_2(mux_tmp_338, mux_tmp_336, nor_tmp_54);
  assign mux_342_nl = MUX_s_1_2_2(mux_tmp_340, mux_340_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_344_nl = MUX_s_1_2_2(mux_tmp_340, mux_342_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_345_nl = MUX_s_1_2_2(mux_tmp_340, mux_344_nl, nor_752_cse);
  assign or_dcpl_147 = mux_345_nl | and_dcpl_779;
  assign or_dcpl_150 = or_dcpl_147 | LOAD_LOOP_for_LOAD_LOOP_nand_cse | and_dcpl_778;
  assign mux_tmp_345 = MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_and_195_ssc_1, or_755_cse,
      or_75_cse);
  assign or_569_nl = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2) | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00)
      | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign nand_37_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 & (~ LOAD_LOOP_for_if_2_for_and_195_ssc_1));
  assign mux_347_nl = MUX_s_1_2_2(or_569_nl, nand_37_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_tmp_419 = LOAD_LOOP_for_if_2_for_or_tmp_1 | mux_347_nl;
  assign mux_tmp_347 = MUX_s_1_2_2(or_tmp_419, or_755_cse, or_75_cse);
  assign mux_tmp_349 = MUX_s_1_2_2(mux_tmp_347, mux_tmp_345, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_349_nl = MUX_s_1_2_2(mux_tmp_347, mux_tmp_345, nor_tmp_54);
  assign mux_351_nl = MUX_s_1_2_2(mux_tmp_349, mux_349_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_353_nl = MUX_s_1_2_2(mux_tmp_349, mux_351_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_tmp_353 = MUX_s_1_2_2(mux_tmp_349, mux_353_nl, nor_752_cse);
  assign or_591_nl = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | LOAD_LOOP_for_if_2_for_equal_tmp_2_1
      | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0]) | (~(or_tmp_154 & (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1])
      & (~ and_tmp_12)));
  assign mux_tmp_359 = MUX_s_1_2_2(or_539_cse, or_591_nl, nor_37_cse);
  assign nand_tmp_41 = ~(and_3266_cse & (~ mux_tmp_359));
  assign or_tmp_471 = nor_566_cse | LOAD_BATCH_LOOP_stage_0 | LOAD_BATCH_LOOP_stage_0_1
      | LOAD_BATCH_LOOP_stage_0_2 | LOAD_BATCH_LOOP_stage_0_3 | (~ LOAD_BATCH_LOOP_stage_v_3);
  assign and_tmp_30 = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1]) & or_tmp_471;
  assign and_tmp_32 = LOAD_LOOP_for_if_2_for_and_195_ssc_1 & or_tmp_471;
  assign nor_tmp_172 = ~(LOAD_BATCH_LOOP_stage_0_1 | (~ LOAD_BATCH_LOOP_stage_v_3));
  assign nor_tmp_175 = or_75_cse & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1]);
  assign mux_tmp_393 = MUX_s_1_2_2(nor_55_cse, (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1]),
      or_75_cse);
  assign mux_tmp_395 = MUX_s_1_2_2(mux_tmp_393, nor_tmp_175, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_395_nl = MUX_s_1_2_2(mux_tmp_393, nor_tmp_175, nor_tmp_54);
  assign mux_397_nl = MUX_s_1_2_2(mux_tmp_395, mux_395_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_399_nl = MUX_s_1_2_2(mux_tmp_395, mux_397_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_tmp_399 = MUX_s_1_2_2(mux_tmp_395, mux_399_nl, nor_752_cse);
  assign or_634_cse = nor_566_cse | LOAD_BATCH_LOOP_stage_0_3 | LOAD_BATCH_LOOP_stage_0_2
      | LOAD_BATCH_LOOP_stage_0;
  assign and_tmp_35 = or_513_cse & or_2860_cse;
  assign or_tmp_497 = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 | (~ or_tmp_471);
  assign nand_279_nl = ~((~((~ LOAD_LOOP_for_asn_6_itm_1) & LOAD_LOOP_for_if_2_for_equal_tmp_1_1))
      & or_tmp_471);
  assign mux_403_nl = MUX_s_1_2_2(or_tmp_497, (~ or_tmp_471), LOAD_LOOP_for_asn_6_itm_1);
  assign mux_404_nl = MUX_s_1_2_2(mux_403_nl, or_tmp_497, dma_read_ctrl_rsci_irdy_mxwt);
  assign mux_405_nl = MUX_s_1_2_2(nand_279_nl, mux_404_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_tmp_405 = MUX_s_1_2_2(mux_405_nl, or_tmp_497, or_750_cse);
  assign not_tmp_236 = ~((lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0==2'b11));
  assign or_682_nl = LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (~(or_tmp_154 & (LOAD_LOOP_for_if_2_for_mux1h_378_tmp==2'b11)
      & (~ and_tmp_12)));
  assign mux_418_nl = MUX_s_1_2_2(or_682_nl, and_tmp_12, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign or_680_nl = exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2
      | not_tmp_236;
  assign mux_tmp_418 = MUX_s_1_2_2(mux_418_nl, or_680_nl, or_75_cse);
  assign nand_tmp_52 = ~(and_3266_cse & (~ mux_tmp_418));
  assign or_tmp_561 = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | LOAD_LOOP_for_LOAD_LOOP_nand_cse;
  assign or_tmp_562 = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | LOAD_LOOP_for_LOAD_LOOP_nand_cse;
  assign mux_tmp_448 = MUX_s_1_2_2(or_tmp_562, or_tmp_561, or_75_cse);
  assign or_731_nl = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2) | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00)
      | or_tmp_562;
  assign nand_58_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 & (~ or_tmp_562));
  assign mux_450_nl = MUX_s_1_2_2(or_731_nl, nand_58_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_tmp_566 = LOAD_LOOP_for_if_2_for_or_tmp_1 | mux_450_nl;
  assign mux_tmp_450 = MUX_s_1_2_2(or_tmp_566, or_tmp_561, or_75_cse);
  assign mux_tmp_452 = MUX_s_1_2_2(mux_tmp_450, mux_tmp_448, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_452_nl = MUX_s_1_2_2(mux_tmp_450, mux_tmp_448, nor_tmp_54);
  assign mux_454_nl = MUX_s_1_2_2(mux_tmp_452, mux_452_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_456_nl = MUX_s_1_2_2(mux_tmp_452, mux_454_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_tmp_456 = MUX_s_1_2_2(mux_tmp_452, mux_456_nl, nor_752_cse);
  assign and_878_nl = or_634_cse & mux_tmp_456;
  assign mux_tmp_457 = MUX_s_1_2_2(mux_tmp_456, and_878_nl, nor_tmp_172);
  assign not_tmp_249 = ~(and_3266_cse & and_tmp_35);
  assign or_tmp_574 = nor_32_cse | (~(LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_nor_tmp
      | (LOAD_BATCH_LOOP_acc_tmp[4]))) | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2)
      | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2
      | not_tmp_249;
  assign nand_tmp_59 = ~(LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse & (~(LOAD_LOOP_for_if_2_for_and_195_ssc_1
      | not_tmp_249)));
  assign or_tmp_577 = nor_32_cse | nand_tmp_59;
  assign mux_tmp_458 = MUX_s_1_2_2(or_tmp_577, or_tmp_574, or_75_cse);
  assign nand_61_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2 & (~(nor_32_cse
      | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00) | nand_tmp_59)));
  assign nand_60_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 & (~ or_tmp_577));
  assign mux_460_nl = MUX_s_1_2_2(nand_61_nl, nand_60_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_747_nl = LOAD_LOOP_for_if_2_for_or_tmp_1 | mux_460_nl;
  assign mux_tmp_460 = MUX_s_1_2_2(or_747_nl, or_tmp_574, or_75_cse);
  assign mux_tmp_462 = MUX_s_1_2_2(mux_tmp_460, mux_tmp_458, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_462_nl = MUX_s_1_2_2(mux_tmp_460, mux_tmp_458, nor_tmp_54);
  assign mux_464_nl = MUX_s_1_2_2(mux_tmp_462, mux_462_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_466_nl = MUX_s_1_2_2(mux_tmp_462, mux_464_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_467_nl = MUX_s_1_2_2(mux_tmp_462, mux_466_nl, nor_752_cse);
  assign nand_tmp_62 = ~(exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0 & (~ mux_467_nl));
  assign mux_tmp_481 = MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_and_195_ssc_1, or_755_cse,
      LOAD_BATCH_LOOP_asn_itm_1);
  assign or_774_nl = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | and_tmp_35;
  assign mux_483_nl = MUX_s_1_2_2(or_755_cse, or_774_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_tmp_483 = MUX_s_1_2_2(mux_483_nl, or_755_cse, nor_32_cse);
  assign mux_tmp_484 = MUX_s_1_2_2(mux_tmp_483, mux_tmp_481, LOAD_BATCH_LOOP_and_3_tmp);
  assign mux_tmp_485 = MUX_s_1_2_2(or_tmp_419, or_755_cse, LOAD_BATCH_LOOP_asn_itm_1);
  assign mux_tmp_486 = MUX_s_1_2_2(mux_tmp_483, mux_tmp_485, LOAD_BATCH_LOOP_and_3_tmp);
  assign nand_tmp_65 = ~(LOAD_BATCH_LOOP_and_3_tmp & (~ mux_tmp_481));
  assign nand_tmp_66 = ~(LOAD_BATCH_LOOP_and_3_tmp & (~ mux_tmp_485));
  assign or_777_nl = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | and_tmp_35;
  assign mux_1158_itm = MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_and_195_ssc_1, or_777_nl,
      LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_tmp_501 = MUX_s_1_2_2(mux_1158_itm, LOAD_LOOP_for_if_2_for_and_195_ssc_1,
      nor_32_cse);
  assign mux_tmp_502 = MUX_s_1_2_2(mux_tmp_501, mux_tmp_483, or_75_cse);
  assign or_tmp_604 = (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00) | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign or_782_nl = (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00) | mux_1158_itm;
  assign mux_504_nl = MUX_s_1_2_2(or_782_nl, or_tmp_604, nor_32_cse);
  assign nand_68_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2 & (~ mux_504_nl));
  assign nand_67_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 & (~ mux_tmp_501));
  assign mux_505_nl = MUX_s_1_2_2(nand_68_nl, nand_67_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_783_nl = LOAD_LOOP_for_if_2_for_or_tmp_1 | mux_505_nl;
  assign mux_tmp_505 = MUX_s_1_2_2(or_783_nl, mux_tmp_483, or_75_cse);
  assign nand_tmp_70 = ~(exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0 & (~ mux_tmp_456));
  assign mux_516_nl = MUX_s_1_2_2(or_tmp_562, or_tmp_561, LOAD_BATCH_LOOP_asn_itm_1);
  assign and_tmp_51 = LOAD_BATCH_LOOP_and_3_tmp & mux_516_nl;
  assign mux_517_nl = MUX_s_1_2_2(or_tmp_566, or_tmp_561, LOAD_BATCH_LOOP_asn_itm_1);
  assign and_tmp_52 = LOAD_BATCH_LOOP_and_3_tmp & mux_517_nl;
  assign mux_tmp_518 = MUX_s_1_2_2(and_tmp_52, and_tmp_51, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_518_nl = MUX_s_1_2_2(and_tmp_52, and_tmp_51, nor_tmp_54);
  assign mux_520_nl = MUX_s_1_2_2(mux_tmp_518, mux_518_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_522_nl = MUX_s_1_2_2(mux_tmp_518, mux_520_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_tmp_522 = MUX_s_1_2_2(mux_tmp_518, mux_522_nl, nor_752_cse);
  assign or_843_cse = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 | LOAD_LOOP_for_if_2_for_equal_tmp_2_1
      | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b10) | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign or_845_nl = nor_tmp_54 | LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b10)
      | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign mux_573_nl = MUX_s_1_2_2(or_843_cse, or_845_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_574_nl = MUX_s_1_2_2(or_843_cse, mux_573_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_575_cse = MUX_s_1_2_2(mux_574_nl, or_843_cse, or_750_cse);
  assign nand_79_nl = ~(or_tmp_154 & (~ mux_575_cse));
  assign mux_tmp_575 = MUX_s_1_2_2(or_539_cse, nand_79_nl, nor_37_cse);
  assign or_872_nl = (~ sfi_operator_8_false_operator_8_false_nor_cse_lpi_2) | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2
      | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b11) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign nand_347_nl = ~(exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_1 & LOAD_LOOP_for_if_2_for_equal_tmp_1
      & LOAD_LOOP_for_if_2_for_mux_11_itm_1 & (~ LOAD_LOOP_for_if_2_for_equal_tmp_1_1));
  assign or_183_nl = (~ LOAD_LOOP_for_if_2_for_mux_11_itm_1) | LOAD_LOOP_for_if_2_for_equal_tmp_1_1;
  assign mux_581_nl = MUX_s_1_2_2(nand_347_nl, or_183_nl, and_3195_cse);
  assign mux_tmp_581 = MUX_s_1_2_2(or_872_nl, mux_581_nl, nor_37_cse);
  assign not_tmp_280 = ~(LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign or_tmp_695 = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | not_tmp_280;
  assign nand_83_nl = ~((~ LOAD_LOOP_for_asn_6_itm_1) & LOAD_LOOP_for_if_2_for_equal_tmp_1_1
      & (~ or_tmp_695));
  assign or_2857_nl = nor_tmp_50 | (~ LOAD_LOOP_for_if_2_for_equal_tmp_1_1) | or_tmp_695;
  assign mux_583_nl = MUX_s_1_2_2(nand_83_nl, or_2857_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign nand_81_nl = ~(LOAD_LOOP_for_if_2_for_equal_tmp_1_1 & (~ or_tmp_695));
  assign mux_tmp_583 = MUX_s_1_2_2(mux_583_nl, nand_81_nl, or_750_cse);
  assign or_tmp_703 = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | (~ and_tmp_35);
  assign or_tmp_704 = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | (~ and_tmp_35);
  assign mux_tmp_589 = MUX_s_1_2_2(or_tmp_704, or_tmp_703, or_75_cse);
  assign or_898_nl = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2) | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00)
      | or_tmp_704;
  assign nand_87_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 & (~ or_tmp_704));
  assign mux_591_nl = MUX_s_1_2_2(or_898_nl, nand_87_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_899_nl = LOAD_LOOP_for_if_2_for_or_tmp_1 | mux_591_nl;
  assign mux_tmp_591 = MUX_s_1_2_2(or_899_nl, or_tmp_703, or_75_cse);
  assign mux_tmp_593 = MUX_s_1_2_2(mux_tmp_591, mux_tmp_589, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_593_nl = MUX_s_1_2_2(mux_tmp_591, mux_tmp_589, nor_tmp_54);
  assign mux_595_nl = MUX_s_1_2_2(mux_tmp_593, mux_593_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_597_nl = MUX_s_1_2_2(mux_tmp_593, mux_595_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_tmp_597 = MUX_s_1_2_2(mux_tmp_593, mux_597_nl, nor_752_cse);
  assign and_dcpl_821 = (~ mux_tmp_597) & LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse
      & or_810_cse;
  assign and_dcpl_831 = and_tmp_25 & LOAD_BATCH_LOOP_stage_v_2 & LOAD_BATCH_LOOP_stage_0_3;
  assign nor_tmp_291 = or_75_cse & exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign or_921_nl = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00)
      | LOAD_LOOP_for_if_2_for_and_195_ssc_1;
  assign mux_603_nl = MUX_s_1_2_2(or_921_nl, or_tmp_151, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_602_nl = MUX_s_1_2_2(or_tmp_604, LOAD_LOOP_for_if_2_for_and_195_ssc_1,
      LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_604_nl = MUX_s_1_2_2(mux_603_nl, mux_602_nl, LOAD_LOOP_for_if_2_for_or_tmp_1);
  assign mux_tmp_604 = MUX_s_1_2_2((~ mux_604_nl), exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2,
      or_75_cse);
  assign nor_695_nl = ~(LOAD_LOOP_if_equal_tmp | (~ or_2860_cse));
  assign or_928_nl = (operator_8_false_7_acc_tmp[8:5]!=4'b0000);
  assign mux_612_itm = MUX_s_1_2_2(nor_695_nl, or_2860_cse, or_928_nl);
  assign or_tmp_723 = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | (~ mux_612_itm);
  assign or_tmp_724 = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | (~ mux_612_itm);
  assign mux_tmp_612 = MUX_s_1_2_2(or_tmp_724, or_tmp_723, or_75_cse);
  assign or_934_nl = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2) | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00)
      | or_tmp_724;
  assign nand_89_nl = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 & (~ or_tmp_724));
  assign mux_614_nl = MUX_s_1_2_2(or_934_nl, nand_89_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_935_nl = LOAD_LOOP_for_if_2_for_or_tmp_1 | mux_614_nl;
  assign mux_tmp_614 = MUX_s_1_2_2(or_935_nl, or_tmp_723, or_75_cse);
  assign or_dcpl_209 = (~ LOAD_LOOP_for_if_2_for_equal_tmp_1) | LOAD_BATCH_LOOP_asn_itm_1
      | (~ LOAD_BATCH_LOOP_and_3_tmp);
  assign or_dcpl_263 = (~(LOAD_LOOP_for_if_2_for_equal_tmp_2_2 & LOAD_BATCH_LOOP_stage_v_2))
      | LOAD_BATCH_LOOP_asn_itm_2 | (~ LOAD_BATCH_LOOP_stage_0_3);
  assign and_tmp_58 = LOAD_LOOP_for_if_2_for_for_and_249_psp & or_tmp_4;
  assign or_tmp_853 = lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2 | (~ exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2)
      | plm_kernel_rsci_bawt;
  assign and_tmp_61 = LOAD_LOOP_for_if_2_for_for_and_248_psp & or_tmp_4;
  assign and_tmp_64 = LOAD_LOOP_for_if_2_for_for_and_247_psp & or_tmp_4;
  assign and_tmp_67 = LOAD_LOOP_for_if_2_for_for_and_246_psp & or_tmp_4;
  assign and_tmp_70 = LOAD_LOOP_for_if_2_for_for_and_245_psp & or_tmp_4;
  assign and_tmp_73 = LOAD_LOOP_for_if_2_for_for_and_244_psp & or_tmp_4;
  assign and_tmp_75 = LOAD_LOOP_for_if_2_for_for_and_243_psp & or_tmp_4;
  assign and_tmp_77 = LOAD_LOOP_for_if_2_for_for_and_242_psp & or_tmp_4;
  assign and_tmp_80 = LOAD_LOOP_for_if_2_for_for_and_241_psp & or_tmp_4;
  assign and_tmp_83 = LOAD_LOOP_for_if_2_for_for_and_240_psp & or_tmp_4;
  assign and_tmp_86 = LOAD_LOOP_for_if_2_for_for_and_239_psp & or_tmp_4;
  assign and_tmp_89 = LOAD_LOOP_for_if_2_for_for_and_238_psp & or_tmp_4;
  assign and_tmp_92 = LOAD_LOOP_for_if_2_for_for_and_237_psp & or_tmp_4;
  assign and_tmp_95 = LOAD_LOOP_for_if_2_for_for_and_236_psp & or_tmp_4;
  assign and_tmp_98 = LOAD_LOOP_for_if_2_for_for_and_235_psp & or_tmp_4;
  assign and_tmp_101 = LOAD_LOOP_for_if_2_for_for_and_234_psp & or_tmp_4;
  assign and_tmp_104 = LOAD_LOOP_for_if_2_for_for_and_233_psp & or_tmp_4;
  assign and_tmp_107 = LOAD_LOOP_for_if_2_for_for_and_232_psp & or_tmp_4;
  assign and_tmp_110 = LOAD_LOOP_for_if_2_for_for_and_231_psp & or_tmp_4;
  assign and_tmp_113 = LOAD_LOOP_for_if_2_for_for_and_230_psp & or_tmp_4;
  assign and_tmp_116 = LOAD_LOOP_for_if_2_for_for_and_229_psp & or_tmp_4;
  assign and_tmp_119 = LOAD_LOOP_for_if_2_for_for_and_228_psp & or_tmp_4;
  assign and_tmp_121 = LOAD_LOOP_for_if_2_for_for_and_227_psp & or_tmp_4;
  assign and_tmp_123 = LOAD_LOOP_for_if_2_for_for_and_226_psp & or_tmp_4;
  assign and_tmp_126 = LOAD_LOOP_for_if_2_for_for_and_225_psp & or_tmp_4;
  assign and_tmp_129 = LOAD_LOOP_for_if_2_for_for_and_224_psp & or_tmp_4;
  assign and_tmp_132 = LOAD_LOOP_for_if_2_for_for_and_223_psp & or_tmp_4;
  assign and_tmp_135 = LOAD_LOOP_for_if_2_for_for_and_222_psp & or_tmp_4;
  assign and_tmp_138 = LOAD_LOOP_for_if_2_for_for_and_221_psp & or_tmp_4;
  assign and_tmp_141 = LOAD_LOOP_for_if_2_for_for_and_220_psp & or_tmp_4;
  assign and_tmp_144 = LOAD_LOOP_for_if_2_for_for_and_219_psp & or_tmp_4;
  assign and_tmp_147 = LOAD_LOOP_for_if_2_for_for_and_218_psp & or_tmp_4;
  assign and_tmp_150 = LOAD_LOOP_for_if_2_for_for_and_217_psp & or_tmp_4;
  assign and_tmp_153 = LOAD_LOOP_for_if_2_for_for_and_216_psp & or_tmp_4;
  assign and_tmp_156 = LOAD_LOOP_for_if_2_for_for_and_215_psp & or_tmp_4;
  assign and_tmp_159 = LOAD_LOOP_for_if_2_for_for_and_214_psp & or_tmp_4;
  assign and_tmp_162 = LOAD_LOOP_for_if_2_for_for_and_213_psp & or_tmp_4;
  assign and_tmp_165 = LOAD_LOOP_for_if_2_for_for_and_212_psp & or_tmp_4;
  assign and_tmp_167 = LOAD_LOOP_for_if_2_for_for_and_211_psp & or_tmp_4;
  assign and_tmp_169 = LOAD_LOOP_for_if_2_for_for_and_210_psp & or_tmp_4;
  assign and_tmp_172 = LOAD_LOOP_for_if_2_for_for_and_209_psp & or_tmp_4;
  assign and_tmp_175 = LOAD_LOOP_for_if_2_for_for_and_208_psp & or_tmp_4;
  assign and_tmp_178 = LOAD_LOOP_for_if_2_for_for_and_207_psp & or_tmp_4;
  assign and_tmp_181 = LOAD_LOOP_for_if_2_for_for_and_206_psp & or_tmp_4;
  assign and_tmp_184 = LOAD_LOOP_for_if_2_for_for_and_205_psp & or_tmp_4;
  assign and_tmp_187 = LOAD_LOOP_for_if_2_for_for_and_204_psp & or_tmp_4;
  assign and_tmp_190 = LOAD_LOOP_for_if_2_for_for_and_203_psp & or_tmp_4;
  assign and_tmp_193 = LOAD_LOOP_for_if_2_for_for_and_202_psp & or_tmp_4;
  assign and_tmp_196 = LOAD_LOOP_for_if_2_for_for_and_201_psp & or_tmp_4;
  assign and_tmp_199 = LOAD_LOOP_for_if_2_for_for_and_200_psp & or_tmp_4;
  assign and_tmp_202 = LOAD_LOOP_for_if_2_for_for_and_199_psp & or_tmp_4;
  assign and_tmp_205 = LOAD_LOOP_for_if_2_for_for_and_198_psp & or_tmp_4;
  assign and_tmp_208 = LOAD_LOOP_for_if_2_for_for_and_197_psp & or_tmp_4;
  assign and_tmp_211 = LOAD_LOOP_for_if_2_for_for_and_196_psp & or_tmp_4;
  assign and_tmp_213 = LOAD_LOOP_for_if_2_for_for_and_195_psp & or_tmp_4;
  assign and_tmp_215 = LOAD_LOOP_for_if_2_for_for_and_194_psp & or_tmp_4;
  assign and_tmp_218 = LOAD_LOOP_for_if_2_for_for_and_193_psp & or_tmp_4;
  assign and_tmp_221 = LOAD_LOOP_for_if_2_for_for_and_192_psp & or_tmp_4;
  assign and_tmp_224 = LOAD_LOOP_for_if_2_for_for_and_191_psp & or_tmp_4;
  assign and_tmp_227 = LOAD_LOOP_for_if_2_for_for_and_190_psp & or_tmp_4;
  assign and_tmp_230 = LOAD_LOOP_for_if_2_for_for_and_189_psp & or_tmp_4;
  assign and_tmp_233 = LOAD_LOOP_for_if_2_for_for_and_188_psp & or_tmp_4;
  assign and_tmp_236 = LOAD_LOOP_for_if_2_for_for_and_187_psp & or_tmp_4;
  assign and_tmp_239 = LOAD_LOOP_for_if_2_for_for_and_186_psp & or_tmp_4;
  assign and_tmp_242 = LOAD_LOOP_for_if_2_for_for_and_185_psp & or_tmp_4;
  assign and_tmp_245 = LOAD_LOOP_for_if_2_for_for_and_184_psp & or_tmp_4;
  assign and_tmp_248 = LOAD_LOOP_for_if_2_for_for_and_183_psp & or_tmp_4;
  assign and_tmp_251 = LOAD_LOOP_for_if_2_for_for_and_182_psp & or_tmp_4;
  assign and_tmp_254 = LOAD_LOOP_for_if_2_for_for_and_181_psp & or_tmp_4;
  assign and_tmp_257 = LOAD_LOOP_for_if_2_for_for_and_180_psp & or_tmp_4;
  assign and_tmp_259 = LOAD_LOOP_for_if_2_for_for_and_179_psp & or_tmp_4;
  assign and_tmp_261 = LOAD_LOOP_for_if_2_for_for_and_178_psp & or_tmp_4;
  assign and_tmp_264 = LOAD_LOOP_for_if_2_for_for_and_177_psp & or_tmp_4;
  assign and_tmp_267 = LOAD_LOOP_for_if_2_for_for_and_176_psp & or_tmp_4;
  assign and_tmp_270 = LOAD_LOOP_for_if_2_for_for_and_175_psp & or_tmp_4;
  assign and_tmp_273 = LOAD_LOOP_for_if_2_for_for_and_174_psp & or_tmp_4;
  assign and_tmp_276 = LOAD_LOOP_for_if_2_for_for_and_173_psp & or_tmp_4;
  assign and_tmp_279 = LOAD_LOOP_for_if_2_for_for_and_172_psp & or_tmp_4;
  assign and_tmp_282 = LOAD_LOOP_for_if_2_for_for_and_171_psp & or_tmp_4;
  assign and_tmp_285 = LOAD_LOOP_for_if_2_for_for_and_170_psp & or_tmp_4;
  assign and_tmp_288 = LOAD_LOOP_for_if_2_for_for_and_169_psp & or_tmp_4;
  assign and_tmp_291 = LOAD_LOOP_for_if_2_for_for_and_168_psp & or_tmp_4;
  assign and_tmp_294 = LOAD_LOOP_for_if_2_for_for_and_167_psp & or_tmp_4;
  assign and_tmp_297 = LOAD_LOOP_for_if_2_for_for_and_166_psp & or_tmp_4;
  assign and_tmp_300 = LOAD_LOOP_for_if_2_for_for_and_165_psp & or_tmp_4;
  assign and_tmp_303 = LOAD_LOOP_for_if_2_for_for_and_164_psp & or_tmp_4;
  assign and_tmp_305 = LOAD_LOOP_for_if_2_for_for_and_163_psp & or_tmp_4;
  assign and_tmp_307 = LOAD_LOOP_for_if_2_for_for_and_162_psp & or_tmp_4;
  assign and_tmp_310 = LOAD_LOOP_for_if_2_for_for_and_161_psp & or_tmp_4;
  assign and_tmp_313 = LOAD_LOOP_for_if_2_for_for_and_160_psp & or_tmp_4;
  assign and_tmp_316 = LOAD_LOOP_for_if_2_for_for_and_159_psp & or_tmp_4;
  assign and_tmp_319 = LOAD_LOOP_for_if_2_for_for_and_158_psp & or_tmp_4;
  assign and_tmp_322 = LOAD_LOOP_for_if_2_for_for_and_157_psp & or_tmp_4;
  assign and_tmp_325 = LOAD_LOOP_for_if_2_for_for_and_156_psp & or_tmp_4;
  assign and_tmp_328 = LOAD_LOOP_for_if_2_for_for_and_155_psp & or_tmp_4;
  assign and_tmp_331 = LOAD_LOOP_for_if_2_for_for_and_154_psp & or_tmp_4;
  assign and_tmp_334 = LOAD_LOOP_for_if_2_for_for_and_153_psp & or_tmp_4;
  assign and_tmp_337 = LOAD_LOOP_for_if_2_for_for_and_152_psp & or_tmp_4;
  assign and_tmp_340 = LOAD_LOOP_for_if_2_for_for_and_151_psp & or_tmp_4;
  assign and_tmp_343 = LOAD_LOOP_for_if_2_for_for_and_150_psp & or_tmp_4;
  assign and_tmp_346 = LOAD_LOOP_for_if_2_for_for_and_149_psp & or_tmp_4;
  assign and_tmp_349 = LOAD_LOOP_for_if_2_for_for_and_148_psp & or_tmp_4;
  assign and_tmp_351 = LOAD_LOOP_for_if_2_for_for_and_147_psp & or_tmp_4;
  assign and_tmp_353 = LOAD_LOOP_for_if_2_for_for_and_146_psp & or_tmp_4;
  assign and_tmp_356 = LOAD_LOOP_for_if_2_for_for_and_145_psp & or_tmp_4;
  assign and_tmp_359 = LOAD_LOOP_for_if_2_for_for_and_144_psp & or_tmp_4;
  assign and_tmp_362 = LOAD_LOOP_for_if_2_for_for_and_143_psp & or_tmp_4;
  assign and_tmp_365 = LOAD_LOOP_for_if_2_for_for_and_142_psp & or_tmp_4;
  assign and_tmp_368 = LOAD_LOOP_for_if_2_for_for_and_141_psp & or_tmp_4;
  assign and_tmp_371 = LOAD_LOOP_for_if_2_for_for_and_140_psp & or_tmp_4;
  assign and_tmp_374 = LOAD_LOOP_for_if_2_for_for_and_139_psp & or_tmp_4;
  assign and_tmp_377 = LOAD_LOOP_for_if_2_for_for_and_138_psp & or_tmp_4;
  assign and_tmp_380 = LOAD_LOOP_for_if_2_for_for_and_137_psp & or_tmp_4;
  assign and_tmp_383 = LOAD_LOOP_for_if_2_for_for_and_136_psp & or_tmp_4;
  assign and_tmp_386 = LOAD_LOOP_for_if_2_for_for_and_135_psp & or_tmp_4;
  assign and_tmp_389 = LOAD_LOOP_for_if_2_for_for_and_134_psp & or_tmp_4;
  assign and_tmp_392 = LOAD_LOOP_for_if_2_for_for_and_133_psp & or_tmp_4;
  assign and_tmp_395 = LOAD_LOOP_for_if_2_for_for_and_132_psp & or_tmp_4;
  assign and_tmp_397 = LOAD_LOOP_for_if_2_for_for_and_131_psp & or_tmp_4;
  assign and_tmp_399 = LOAD_LOOP_for_if_2_for_for_and_130_psp & or_tmp_4;
  assign and_tmp_402 = LOAD_LOOP_for_if_2_for_for_and_129_psp & or_tmp_4;
  assign and_tmp_405 = LOAD_LOOP_for_if_2_for_for_and_128_psp & or_tmp_4;
  assign and_tmp_408 = LOAD_LOOP_for_if_2_for_for_and_127_psp & or_tmp_4;
  assign and_tmp_411 = LOAD_LOOP_for_if_2_for_for_and_126_psp & or_tmp_4;
  assign and_tmp_414 = LOAD_LOOP_for_if_2_for_for_and_125_psp & or_tmp_4;
  assign and_tmp_417 = LOAD_LOOP_for_if_2_for_for_and_124_psp & or_tmp_4;
  assign mux_93_nl = MUX_s_1_2_2(mux_tmp_91, and_tmp_17, nor_tmp_54);
  assign mux_95_nl = MUX_s_1_2_2(mux_tmp_93, mux_93_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_97_nl = MUX_s_1_2_2(mux_tmp_93, mux_95_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_98_nl = MUX_s_1_2_2(mux_tmp_93, mux_97_nl, nor_752_cse);
  assign or_tmp_1480 = (mux_98_nl | LOAD_LOOP_for_LOAD_LOOP_nand_cse) & LOAD_BATCH_LOOP_and_4_tmp
      & (fsm_output[2]);
  assign or_tmp_1481 = (~ mux_tmp_581) & and_dcpl_28 & (fsm_output[2]);
  assign or_439_cse = (~ operator_8_false_operator_8_false_nor_cse_lpi_2) | (~ LOAD_LOOP_for_if_2_for_for_if_aelse_2_acc_itm_9_1)
      | (~ LOAD_LOOP_for_if_2_for_for_if_aelse_1_acc_itm_9_1) | LOAD_LOOP_for_if_2_for_for_if_aelse_acc_itm_8
      | (z_out_11[8]);
  assign or_447_nl = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b10) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign or_446_nl = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign mux_257_nl = MUX_s_1_2_2(or_447_nl, or_446_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2);
  assign mux_253_nl = MUX_s_1_2_2(or_tmp_325, LOAD_LOOP_for_if_2_for_and_195_ssc_1,
      LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1]);
  assign mux_252_nl = MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_and_195_ssc_1, or_tmp_325,
      LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1]);
  assign mux_254_nl = MUX_s_1_2_2(mux_253_nl, mux_252_nl, nor_tmp_67);
  assign mux_255_nl = MUX_s_1_2_2(mux_254_nl, or_tmp_325, LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0]);
  assign mux_251_nl = MUX_s_1_2_2(or_tmp_325, LOAD_LOOP_for_if_2_for_and_195_ssc_1,
      nor_tmp_63);
  assign mux_256_nl = MUX_s_1_2_2(mux_255_nl, mux_251_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_258_nl = MUX_s_1_2_2(mux_257_nl, mux_256_nl, nor_37_cse);
  assign or_443_nl = LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0])
      | (~(nor_113_cse & (~(LOAD_LOOP_for_if_2_for_and_195_ssc_1 | and_tmp_12))));
  assign mux_250_nl = MUX_s_1_2_2(or_539_cse, or_443_nl, nor_37_cse);
  assign mux_259_nl = MUX_s_1_2_2(mux_258_nl, mux_250_nl, or_439_cse);
  assign or_tmp_2017 = (~ mux_259_nl) & and_dcpl_752 & (fsm_output[2]);
  assign nor_778_cse = ~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b10)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2);
  assign or_tmp_2027 = or_tmp_4 & ((~ LOAD_BATCH_LOOP_and_3_tmp) | (~ exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_1)
      | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0]) | or_dcpl_34) &
      and_dcpl_764 & (fsm_output[2]);
  assign or_tmp_2033 = (or_dcpl_122 | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1])
      | (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2 & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_2))
      | and_dcpl_186 | (~(LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_2
      & LOAD_BATCH_LOOP_stage_0_3))) & and_dcpl_772 & (fsm_output[2]);
  assign or_tmp_2041 = (~ (fsm_output[2])) | or_dcpl_129 | (~(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2
      & LOAD_LOOP_for_if_2_for_for_asn_itm_1));
  assign or_588_cse = nor_566_cse | LOAD_BATCH_LOOP_stage_0_1 | (~ LOAD_BATCH_LOOP_stage_v_3)
      | LOAD_BATCH_LOOP_stage_0_3 | LOAD_BATCH_LOOP_stage_0_2;
  assign mux_364_nl = MUX_s_1_2_2((~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1])),
      (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1]), lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2);
  assign or_604_nl = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[0]) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2
      | mux_364_nl;
  assign nand_43_nl = ~((LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1]) & (~ and_tmp_12));
  assign or_601_nl = (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1]) | and_tmp_12;
  assign mux_361_nl = MUX_s_1_2_2(nand_43_nl, or_601_nl, or_tmp_154);
  assign mux_362_nl = MUX_s_1_2_2(mux_361_nl, and_tmp_12, LOAD_LOOP_for_if_2_for_mux1h_378_tmp[0]);
  assign nand_42_nl = ~(or_tmp_388 & (~ and_tmp_12));
  assign mux_363_nl = MUX_s_1_2_2(mux_362_nl, nand_42_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign or_602_nl = LOAD_LOOP_for_if_2_for_and_195_ssc_1 | (~ mux_363_nl);
  assign mux_365_nl = MUX_s_1_2_2(or_604_nl, or_602_nl, nor_37_cse);
  assign mux_366_nl = MUX_s_1_2_2(mux_tmp_359, mux_365_nl, or_2860_cse);
  assign mux_367_nl = MUX_s_1_2_2(mux_tmp_359, mux_366_nl, or_513_cse);
  assign nand_44_nl = ~(and_3266_cse & (~ mux_367_nl));
  assign mux_368_nl = MUX_s_1_2_2(nand_tmp_41, nand_44_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, nand_tmp_41, nor_32_cse);
  assign mux_370_nl = MUX_s_1_2_2(nand_tmp_41, mux_369_nl, exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign and_840_nl = LOAD_BATCH_LOOP_stage_0 & mux_370_nl;
  assign mux_371_nl = MUX_s_1_2_2(and_840_nl, nand_tmp_41, or_588_cse);
  assign or_tmp_2056 = mux_371_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign or_tmp_2094 = mux_tmp_457 & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign and_3252_nl = or_tmp_154 & (~ mux_575_cse);
  assign mux_580_nl = MUX_s_1_2_2(nor_778_cse, and_3252_nl, nor_37_cse);
  assign or_tmp_2314 = mux_580_nl & and_dcpl_752 & (fsm_output[2]);
  assign or_tmp_2315 = (mux_tmp_575 | LOAD_LOOP_for_LOAD_LOOP_nand_cse) & LOAD_BATCH_LOOP_and_4_tmp
      & (fsm_output[2]);
  assign or_tmp_2337 = (~ LOAD_BATCH_LOOP_asn_itm_1) & LOAD_BATCH_LOOP_and_3_tmp
      & (fsm_output[2]);
  assign or_tmp_2350 = and_dcpl_821 & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0
      & and_dcpl_752 & (fsm_output[2]);
  assign or_tmp_2354 = nand_tmp_62 & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign or_189_nl = sfi_operator_8_false_operator_8_false_nor_cse_lpi_2 | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2
      | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b11) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign nand_23_nl = ~(LOAD_LOOP_for_if_2_for_and_195_ssc_1 & (~ mux_tmp_103));
  assign mux_105_nl = MUX_s_1_2_2(nand_23_nl, mux_tmp_103, and_3195_cse);
  assign mux_106_nl = MUX_s_1_2_2(or_189_nl, mux_105_nl, nor_37_cse);
  assign dma_read_ctrl_rsci_idat_15_0_mx0c2 = (~ mux_106_nl) & and_dcpl_28 & (fsm_output[2]);
  assign dma_read_ctrl_rsci_idat_47_32_mx0c1 = (~ mux_481_cse) & and_dcpl_28 & (fsm_output[2]);
  assign plm_kernel_rsci_idat_31_0_mx0c1 = (or_dcpl_32 | or_dcpl_30) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_63_32_mx0c1 = (or_dcpl_32 | or_dcpl_39) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_95_64_mx0c1 = (or_dcpl_32 | or_dcpl_42) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_127_96_mx0c1 = (or_dcpl_32 | or_dcpl_45) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_159_128_mx0c1 = (or_dcpl_32 | or_dcpl_47) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_191_160_mx0c1 = (or_dcpl_32 | or_dcpl_49) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_223_192_mx0c1 = (or_dcpl_32 | or_dcpl_51) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_255_224_mx0c1 = (or_dcpl_32 | or_dcpl_53) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_287_256_mx0c1 = (or_dcpl_56 | or_dcpl_30) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_319_288_mx0c1 = (or_dcpl_56 | or_dcpl_39) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_351_320_mx0c1 = (or_dcpl_56 | or_dcpl_42) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_383_352_mx0c1 = (or_dcpl_56 | or_dcpl_45) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_415_384_mx0c1 = (or_dcpl_56 | or_dcpl_47) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_447_416_mx0c1 = (or_dcpl_56 | or_dcpl_49) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_479_448_mx0c1 = (or_dcpl_56 | or_dcpl_51) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_511_480_mx0c1 = (or_dcpl_56 | or_dcpl_53) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_543_512_mx0c1 = (or_dcpl_66 | or_dcpl_30) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_575_544_mx0c1 = (or_dcpl_66 | or_dcpl_39) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_607_576_mx0c1 = (or_dcpl_66 | or_dcpl_42) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_639_608_mx0c1 = (or_dcpl_66 | or_dcpl_45) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_671_640_mx0c1 = (or_dcpl_66 | or_dcpl_47) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_703_672_mx0c1 = (or_dcpl_66 | or_dcpl_49) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_735_704_mx0c1 = (or_dcpl_66 | or_dcpl_51) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_767_736_mx0c1 = (or_dcpl_66 | or_dcpl_53) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_799_768_mx0c1 = (or_dcpl_76 | or_dcpl_30) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_831_800_mx0c1 = (or_dcpl_76 | or_dcpl_39) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_863_832_mx0c1 = (or_dcpl_76 | or_dcpl_42) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_895_864_mx0c1 = (or_dcpl_76 | or_dcpl_45) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_927_896_mx0c1 = (or_dcpl_76 | or_dcpl_47) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_959_928_mx0c1 = (or_dcpl_76 | or_dcpl_49) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_991_960_mx0c1 = (or_dcpl_76 | or_dcpl_51) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1023_992_mx0c1 = (or_dcpl_76 | or_dcpl_53) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1055_1024_mx0c1 = (or_dcpl_85 | or_dcpl_30) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1087_1056_mx0c1 = (or_dcpl_85 | or_dcpl_39) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1119_1088_mx0c1 = (or_dcpl_85 | or_dcpl_42) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1151_1120_mx0c1 = (or_dcpl_85 | or_dcpl_45) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1183_1152_mx0c1 = (or_dcpl_85 | or_dcpl_47) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1215_1184_mx0c1 = (or_dcpl_85 | or_dcpl_49) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1247_1216_mx0c1 = (or_dcpl_85 | or_dcpl_51) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1279_1248_mx0c1 = (or_dcpl_85 | or_dcpl_53) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1311_1280_mx0c1 = (or_dcpl_94 | or_dcpl_30) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1343_1312_mx0c1 = (or_dcpl_94 | or_dcpl_39) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1375_1344_mx0c1 = (or_dcpl_94 | or_dcpl_42) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1407_1376_mx0c1 = (or_dcpl_94 | or_dcpl_45) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1439_1408_mx0c1 = (or_dcpl_94 | or_dcpl_47) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1471_1440_mx0c1 = (or_dcpl_94 | or_dcpl_49) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1503_1472_mx0c1 = (or_dcpl_94 | or_dcpl_51) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1535_1504_mx0c1 = (or_dcpl_94 | or_dcpl_53) & and_dcpl_44
      & (fsm_output[2]);
  assign plm_kernel_rsci_idat_1567_1536_mx0c1 = (or_dcpl_103 | or_dcpl_30) & and_dcpl_44
      & (fsm_output[2]);
  assign or_289_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000);
  assign mux_124_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_289_cse);
  assign buf_linear_rsci_idat_31_0_mx0c1 = mux_124_nl & or_9_cse & and_dcpl_183 &
      (fsm_output[2]);
  assign mux_125_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_289_cse);
  assign buf_linear_rsci_idat_63_32_mx0c1 = mux_125_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_126_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_289_cse);
  assign buf_linear_rsci_idat_95_64_mx0c1 = mux_126_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_127_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_289_cse);
  assign buf_linear_rsci_idat_127_96_mx0c1 = mux_127_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_305_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000);
  assign mux_128_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_305_cse);
  assign buf_linear_rsci_idat_159_128_mx0c1 = mux_128_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_129_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_305_cse);
  assign buf_linear_rsci_idat_191_160_mx0c1 = mux_129_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_130_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_305_cse);
  assign buf_linear_rsci_idat_223_192_mx0c1 = mux_130_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_131_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_305_cse);
  assign buf_linear_rsci_idat_255_224_mx0c1 = mux_131_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_309_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000);
  assign mux_132_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_309_cse);
  assign buf_linear_rsci_idat_287_256_mx0c1 = mux_132_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_133_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_309_cse);
  assign buf_linear_rsci_idat_319_288_mx0c1 = mux_133_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_134_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_309_cse);
  assign buf_linear_rsci_idat_351_320_mx0c1 = mux_134_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_135_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_309_cse);
  assign buf_linear_rsci_idat_383_352_mx0c1 = mux_135_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_313_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b11)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000);
  assign mux_136_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_313_cse);
  assign buf_linear_rsci_idat_415_384_mx0c1 = mux_136_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_137_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_313_cse);
  assign buf_linear_rsci_idat_447_416_mx0c1 = mux_137_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_138_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_313_cse);
  assign buf_linear_rsci_idat_479_448_mx0c1 = mux_138_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_139_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_313_cse);
  assign buf_linear_rsci_idat_511_480_mx0c1 = mux_139_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_317_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001);
  assign mux_140_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_317_cse);
  assign buf_linear_rsci_idat_543_512_mx0c1 = mux_140_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_141_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_317_cse);
  assign buf_linear_rsci_idat_575_544_mx0c1 = mux_141_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_142_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_317_cse);
  assign buf_linear_rsci_idat_607_576_mx0c1 = mux_142_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_143_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_317_cse);
  assign buf_linear_rsci_idat_639_608_mx0c1 = mux_143_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_321_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001);
  assign mux_144_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_321_cse);
  assign buf_linear_rsci_idat_671_640_mx0c1 = mux_144_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_145_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_321_cse);
  assign buf_linear_rsci_idat_703_672_mx0c1 = mux_145_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_146_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_321_cse);
  assign buf_linear_rsci_idat_735_704_mx0c1 = mux_146_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_147_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_321_cse);
  assign buf_linear_rsci_idat_767_736_mx0c1 = mux_147_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_325_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001);
  assign mux_148_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_325_cse);
  assign buf_linear_rsci_idat_799_768_mx0c1 = mux_148_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_149_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_325_cse);
  assign buf_linear_rsci_idat_831_800_mx0c1 = mux_149_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_150_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_325_cse);
  assign buf_linear_rsci_idat_863_832_mx0c1 = mux_150_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_151_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_325_cse);
  assign buf_linear_rsci_idat_895_864_mx0c1 = mux_151_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_329_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b11)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001);
  assign mux_152_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_329_cse);
  assign buf_linear_rsci_idat_927_896_mx0c1 = mux_152_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_153_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_329_cse);
  assign buf_linear_rsci_idat_959_928_mx0c1 = mux_153_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_154_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_329_cse);
  assign buf_linear_rsci_idat_991_960_mx0c1 = mux_154_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_155_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_329_cse);
  assign buf_linear_rsci_idat_1023_992_mx0c1 = mux_155_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_333_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010);
  assign mux_156_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_333_cse);
  assign buf_linear_rsci_idat_1055_1024_mx0c1 = mux_156_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_157_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_333_cse);
  assign buf_linear_rsci_idat_1087_1056_mx0c1 = mux_157_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_158_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_333_cse);
  assign buf_linear_rsci_idat_1119_1088_mx0c1 = mux_158_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_159_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_333_cse);
  assign buf_linear_rsci_idat_1151_1120_mx0c1 = mux_159_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_337_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010);
  assign mux_160_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_337_cse);
  assign buf_linear_rsci_idat_1183_1152_mx0c1 = mux_160_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_161_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_337_cse);
  assign buf_linear_rsci_idat_1215_1184_mx0c1 = mux_161_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_162_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_337_cse);
  assign buf_linear_rsci_idat_1247_1216_mx0c1 = mux_162_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_163_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_337_cse);
  assign buf_linear_rsci_idat_1279_1248_mx0c1 = mux_163_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_341_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010);
  assign mux_164_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_341_cse);
  assign buf_linear_rsci_idat_1311_1280_mx0c1 = mux_164_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_165_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_341_cse);
  assign buf_linear_rsci_idat_1343_1312_mx0c1 = mux_165_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_166_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_341_cse);
  assign buf_linear_rsci_idat_1375_1344_mx0c1 = mux_166_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_167_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_341_cse);
  assign buf_linear_rsci_idat_1407_1376_mx0c1 = mux_167_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_345_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b11)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010);
  assign mux_168_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_345_cse);
  assign buf_linear_rsci_idat_1439_1408_mx0c1 = mux_168_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_169_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_345_cse);
  assign buf_linear_rsci_idat_1471_1440_mx0c1 = mux_169_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_170_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_345_cse);
  assign buf_linear_rsci_idat_1503_1472_mx0c1 = mux_170_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_171_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_345_cse);
  assign buf_linear_rsci_idat_1535_1504_mx0c1 = mux_171_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_349_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011);
  assign mux_172_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_349_cse);
  assign buf_linear_rsci_idat_1567_1536_mx0c1 = mux_172_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_173_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_349_cse);
  assign buf_linear_rsci_idat_1599_1568_mx0c1 = mux_173_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_174_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_349_cse);
  assign buf_linear_rsci_idat_1631_1600_mx0c1 = mux_174_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_175_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_349_cse);
  assign buf_linear_rsci_idat_1663_1632_mx0c1 = mux_175_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_353_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011);
  assign mux_176_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_353_cse);
  assign buf_linear_rsci_idat_1695_1664_mx0c1 = mux_176_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_177_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_353_cse);
  assign buf_linear_rsci_idat_1727_1696_mx0c1 = mux_177_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_178_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_353_cse);
  assign buf_linear_rsci_idat_1759_1728_mx0c1 = mux_178_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_179_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_353_cse);
  assign buf_linear_rsci_idat_1791_1760_mx0c1 = mux_179_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_357_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011);
  assign mux_180_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, or_357_cse);
  assign buf_linear_rsci_idat_1823_1792_mx0c1 = mux_180_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_181_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, or_357_cse);
  assign buf_linear_rsci_idat_1855_1824_mx0c1 = mux_181_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_182_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, or_357_cse);
  assign buf_linear_rsci_idat_1887_1856_mx0c1 = mux_182_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_183_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, or_357_cse);
  assign buf_linear_rsci_idat_1919_1888_mx0c1 = mux_183_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign nand_106_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b011));
  assign mux_184_nl = MUX_s_1_2_2(not_tmp_118, or_tmp_4, nand_106_cse);
  assign buf_linear_rsci_idat_1951_1920_mx0c1 = mux_184_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_185_nl = MUX_s_1_2_2(not_tmp_124, or_tmp_4, nand_106_cse);
  assign buf_linear_rsci_idat_1983_1952_mx0c1 = mux_185_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_186_nl = MUX_s_1_2_2(not_tmp_125, or_tmp_4, nand_106_cse);
  assign buf_linear_rsci_idat_2015_1984_mx0c1 = mux_186_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_187_nl = MUX_s_1_2_2(not_tmp_126, or_tmp_4, nand_106_cse);
  assign buf_linear_rsci_idat_2047_2016_mx0c1 = mux_187_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_365_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]!=2'b00);
  assign mux_188_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, or_365_cse);
  assign buf_linear_rsci_idat_2079_2048_mx0c1 = mux_188_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_189_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, or_365_cse);
  assign buf_linear_rsci_idat_2111_2080_mx0c1 = mux_189_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_190_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, or_365_cse);
  assign buf_linear_rsci_idat_2143_2112_mx0c1 = mux_190_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_191_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, or_365_cse);
  assign buf_linear_rsci_idat_2175_2144_mx0c1 = mux_191_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_373_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]!=2'b00);
  assign mux_192_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, or_373_cse);
  assign buf_linear_rsci_idat_2207_2176_mx0c1 = mux_192_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_193_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, or_373_cse);
  assign buf_linear_rsci_idat_2239_2208_mx0c1 = mux_193_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_194_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, or_373_cse);
  assign buf_linear_rsci_idat_2271_2240_mx0c1 = mux_194_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_195_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, or_373_cse);
  assign buf_linear_rsci_idat_2303_2272_mx0c1 = mux_195_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_377_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]!=2'b00);
  assign mux_196_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, or_377_cse);
  assign buf_linear_rsci_idat_2335_2304_mx0c1 = mux_196_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_197_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, or_377_cse);
  assign buf_linear_rsci_idat_2367_2336_mx0c1 = mux_197_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_198_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, or_377_cse);
  assign buf_linear_rsci_idat_2399_2368_mx0c1 = mux_198_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_199_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, or_377_cse);
  assign buf_linear_rsci_idat_2431_2400_mx0c1 = mux_199_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_381_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b11)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]!=2'b00);
  assign mux_200_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, or_381_cse);
  assign buf_linear_rsci_idat_2463_2432_mx0c1 = mux_200_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_201_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, or_381_cse);
  assign buf_linear_rsci_idat_2495_2464_mx0c1 = mux_201_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_202_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, or_381_cse);
  assign buf_linear_rsci_idat_2527_2496_mx0c1 = mux_202_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_203_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, or_381_cse);
  assign buf_linear_rsci_idat_2559_2528_mx0c1 = mux_203_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_385_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]!=2'b01);
  assign mux_204_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, or_385_cse);
  assign buf_linear_rsci_idat_2591_2560_mx0c1 = mux_204_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_205_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, or_385_cse);
  assign buf_linear_rsci_idat_2623_2592_mx0c1 = mux_205_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_206_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, or_385_cse);
  assign buf_linear_rsci_idat_2655_2624_mx0c1 = mux_206_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_207_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, or_385_cse);
  assign buf_linear_rsci_idat_2687_2656_mx0c1 = mux_207_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_389_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]!=2'b01);
  assign mux_208_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, or_389_cse);
  assign buf_linear_rsci_idat_2719_2688_mx0c1 = mux_208_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_209_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, or_389_cse);
  assign buf_linear_rsci_idat_2751_2720_mx0c1 = mux_209_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_210_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, or_389_cse);
  assign buf_linear_rsci_idat_2783_2752_mx0c1 = mux_210_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_211_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, or_389_cse);
  assign buf_linear_rsci_idat_2815_2784_mx0c1 = mux_211_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_393_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]!=2'b01);
  assign mux_212_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, or_393_cse);
  assign buf_linear_rsci_idat_2847_2816_mx0c1 = mux_212_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_213_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, or_393_cse);
  assign buf_linear_rsci_idat_2879_2848_mx0c1 = mux_213_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_214_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, or_393_cse);
  assign buf_linear_rsci_idat_2911_2880_mx0c1 = mux_214_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_215_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, or_393_cse);
  assign buf_linear_rsci_idat_2943_2912_mx0c1 = mux_215_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign nand_102_cse = ~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]==2'b01));
  assign mux_216_nl = MUX_s_1_2_2(not_tmp_127, or_tmp_4, nand_102_cse);
  assign buf_linear_rsci_idat_2975_2944_mx0c1 = mux_216_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_217_nl = MUX_s_1_2_2(not_tmp_128, or_tmp_4, nand_102_cse);
  assign buf_linear_rsci_idat_3007_2976_mx0c1 = mux_217_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_218_nl = MUX_s_1_2_2(not_tmp_129, or_tmp_4, nand_102_cse);
  assign buf_linear_rsci_idat_3039_3008_mx0c1 = mux_218_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_219_nl = MUX_s_1_2_2(not_tmp_130, or_tmp_4, nand_102_cse);
  assign buf_linear_rsci_idat_3071_3040_mx0c1 = mux_219_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_401_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign mux_220_nl = MUX_s_1_2_2(not_tmp_131, or_tmp_4, or_401_cse);
  assign buf_linear_rsci_idat_3103_3072_mx0c1 = mux_220_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_221_nl = MUX_s_1_2_2(not_tmp_132, or_tmp_4, or_401_cse);
  assign buf_linear_rsci_idat_3135_3104_mx0c1 = mux_221_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_222_nl = MUX_s_1_2_2(not_tmp_133, or_tmp_4, or_401_cse);
  assign buf_linear_rsci_idat_3167_3136_mx0c1 = mux_222_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_223_nl = MUX_s_1_2_2(not_tmp_134, or_tmp_4, or_401_cse);
  assign buf_linear_rsci_idat_3199_3168_mx0c1 = mux_223_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_409_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign mux_224_nl = MUX_s_1_2_2(not_tmp_131, or_tmp_4, or_409_cse);
  assign buf_linear_rsci_idat_3231_3200_mx0c1 = mux_224_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_225_nl = MUX_s_1_2_2(not_tmp_132, or_tmp_4, or_409_cse);
  assign buf_linear_rsci_idat_3263_3232_mx0c1 = mux_225_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_226_nl = MUX_s_1_2_2(not_tmp_133, or_tmp_4, or_409_cse);
  assign buf_linear_rsci_idat_3295_3264_mx0c1 = mux_226_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_227_nl = MUX_s_1_2_2(not_tmp_134, or_tmp_4, or_409_cse);
  assign buf_linear_rsci_idat_3327_3296_mx0c1 = mux_227_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_413_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign mux_228_nl = MUX_s_1_2_2(not_tmp_131, or_tmp_4, or_413_cse);
  assign buf_linear_rsci_idat_3359_3328_mx0c1 = mux_228_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_229_nl = MUX_s_1_2_2(not_tmp_132, or_tmp_4, or_413_cse);
  assign buf_linear_rsci_idat_3391_3360_mx0c1 = mux_229_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_230_nl = MUX_s_1_2_2(not_tmp_133, or_tmp_4, or_413_cse);
  assign buf_linear_rsci_idat_3423_3392_mx0c1 = mux_230_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_231_nl = MUX_s_1_2_2(not_tmp_134, or_tmp_4, or_413_cse);
  assign buf_linear_rsci_idat_3455_3424_mx0c1 = mux_231_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_417_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b11)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[0]);
  assign mux_232_nl = MUX_s_1_2_2(not_tmp_131, or_tmp_4, or_417_cse);
  assign buf_linear_rsci_idat_3487_3456_mx0c1 = mux_232_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_233_nl = MUX_s_1_2_2(not_tmp_132, or_tmp_4, or_417_cse);
  assign buf_linear_rsci_idat_3519_3488_mx0c1 = mux_233_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_234_nl = MUX_s_1_2_2(not_tmp_133, or_tmp_4, or_417_cse);
  assign buf_linear_rsci_idat_3551_3520_mx0c1 = mux_234_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_235_nl = MUX_s_1_2_2(not_tmp_134, or_tmp_4, or_417_cse);
  assign buf_linear_rsci_idat_3583_3552_mx0c1 = mux_235_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_421_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00);
  assign mux_236_nl = MUX_s_1_2_2(not_tmp_135, or_tmp_4, or_421_cse);
  assign buf_linear_rsci_idat_3615_3584_mx0c1 = mux_236_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_237_nl = MUX_s_1_2_2(not_tmp_136, or_tmp_4, or_421_cse);
  assign buf_linear_rsci_idat_3647_3616_mx0c1 = mux_237_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_238_nl = MUX_s_1_2_2(not_tmp_137, or_tmp_4, or_421_cse);
  assign buf_linear_rsci_idat_3679_3648_mx0c1 = mux_238_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_239_nl = MUX_s_1_2_2(not_tmp_138, or_tmp_4, or_421_cse);
  assign buf_linear_rsci_idat_3711_3680_mx0c1 = mux_239_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign or_429_cse = (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b01);
  assign mux_240_nl = MUX_s_1_2_2(not_tmp_135, or_tmp_4, or_429_cse);
  assign buf_linear_rsci_idat_3743_3712_mx0c1 = mux_240_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_241_nl = MUX_s_1_2_2(not_tmp_136, or_tmp_4, or_429_cse);
  assign buf_linear_rsci_idat_3775_3744_mx0c1 = mux_241_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_242_nl = MUX_s_1_2_2(not_tmp_137, or_tmp_4, or_429_cse);
  assign buf_linear_rsci_idat_3807_3776_mx0c1 = mux_242_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign mux_243_nl = MUX_s_1_2_2(not_tmp_138, or_tmp_4, or_429_cse);
  assign buf_linear_rsci_idat_3839_3808_mx0c1 = mux_243_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign and_3202_nl = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1)) & or_tmp_4;
  assign mux_244_nl = MUX_s_1_2_2(and_3202_nl, or_tmp_4, LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign buf_linear_rsci_idat_3871_3840_mx0c1 = mux_244_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign and_3201_nl = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1)) & or_tmp_4;
  assign mux_245_nl = MUX_s_1_2_2(and_3201_nl, or_tmp_4, LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign buf_linear_rsci_idat_3903_3872_mx0c1 = mux_245_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign and_3200_nl = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1)) & or_tmp_4;
  assign mux_246_nl = MUX_s_1_2_2(and_3200_nl, or_tmp_4, LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign buf_linear_rsci_idat_3935_3904_mx0c1 = mux_246_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign and_3199_nl = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1)) & or_tmp_4;
  assign mux_247_nl = MUX_s_1_2_2(and_3199_nl, or_tmp_4, LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]);
  assign buf_linear_rsci_idat_3967_3936_mx0c1 = mux_247_nl & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign buf_linear_rsci_idat_3999_3968_mx0c1 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1)) & or_tmp_4 & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign buf_linear_rsci_idat_4031_4000_mx0c1 = (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1)) & or_tmp_4 & or_9_cse & and_dcpl_183
      & (fsm_output[2]);
  assign and_893_nl = LOAD_BATCH_LOOP_stage_0 & nand_tmp_70;
  assign mux_524_nl = MUX_s_1_2_2(LOAD_BATCH_LOOP_and_3_tmp, mux_tmp_522, exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign mux_525_nl = MUX_s_1_2_2(mux_524_nl, nand_tmp_70, LOAD_BATCH_LOOP_stage_0);
  assign mux_526_nl = MUX_s_1_2_2(and_893_nl, mux_525_nl, LOAD_BATCH_LOOP_stage_0_2);
  assign mux_527_nl = MUX_s_1_2_2(mux_526_nl, nand_tmp_70, or_771_cse);
  assign mux_528_nl = MUX_s_1_2_2(mux_527_nl, nand_tmp_70, LOAD_BATCH_LOOP_stage_0_1);
  assign LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1_mx0c1 = mux_528_nl
      & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2_mx0c1 = (mux_tmp_581 | LOAD_LOOP_for_LOAD_LOOP_nand_cse
      | (~ LOAD_LOOP_for_asn_sft_lpi_2)) & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign or_889_nl = (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00)
      | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | not_tmp_280;
  assign mux_586_nl = MUX_s_1_2_2(or_tmp_695, mux_tmp_583, or_101_cse);
  assign mux_585_nl = MUX_s_1_2_2(or_tmp_695, mux_tmp_583, or_93_cse);
  assign mux_587_nl = MUX_s_1_2_2(mux_586_nl, mux_585_nl, or_44_cse);
  assign mux_588_nl = MUX_s_1_2_2(or_889_nl, mux_587_nl, nor_37_cse);
  assign nand_86_nl = ~(or_810_cse & or_513_cse & or_2860_cse & lfst_exit_LOAD_LOOP_for_1_lpi_2
      & lfst_exit_LOAD_LOOP_sva & (~ mux_588_nl));
  assign mux_589_nl = MUX_s_1_2_2((~ LOAD_BATCH_LOOP_stage_v), nand_86_nl, LOAD_BATCH_LOOP_and_4_tmp);
  assign LOAD_BATCH_LOOP_stage_v_mx0c0 = (fsm_output[1]) | (mux_589_nl & LOAD_BATCH_LOOP_stage_0
      & (fsm_output[2]));
  assign LOAD_BATCH_LOOP_stage_v_mx0c1 = (~((~(and_dcpl_821 & and_3266_cse & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0))
      & LOAD_BATCH_LOOP_stage_0)) & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign LOAD_BATCH_LOOP_stage_v_2_mx0c0 = (fsm_output[1]) | (and_tmp_25 & LOAD_BATCH_LOOP_stage_v_2
      & (~ LOAD_BATCH_LOOP_and_3_tmp) & LOAD_BATCH_LOOP_stage_0_3 & (fsm_output[2]));
  assign and_3222_nl = or_42_cse & LOAD_BATCH_LOOP_stage_v_2;
  assign and_3223_nl = or_41_cse & LOAD_BATCH_LOOP_stage_v_2;
  assign mux_599_nl = MUX_s_1_2_2(and_3222_nl, and_3223_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_3224_nl = or_tmp_57 & LOAD_BATCH_LOOP_stage_v_2;
  assign mux_600_nl = MUX_s_1_2_2(mux_599_nl, and_3224_nl, or_9_cse);
  assign LOAD_BATCH_LOOP_stage_v_3_mx0c0 = (fsm_output[1]) | ((~(nor_566_cse | (LOAD_BATCH_LOOP_stage_0_3
      & mux_600_nl))) & LOAD_BATCH_LOOP_stage_v_3 & (fsm_output[2]));
  assign LOAD_LOOP_for_k_5_0_lpi_2_4_0_mx0c1 = or_dcpl_150 & LOAD_BATCH_LOOP_and_4_tmp;
  assign LOAD_BATCH_LOOP_stage_v_1_mx0c0 = (fsm_output[1]) | (LOAD_BATCH_LOOP_and_3_tmp
      & (~ LOAD_BATCH_LOOP_and_4_tmp) & (fsm_output[2]));
  assign nl_LOAD_LOOP_for_if_2_for_for_if_aelse_acc_nl = ({4'b1000 , LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1})
      + conv_u2u_8_9(~ pad_sva) + 9'b000000001;
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_acc_nl = nl_LOAD_LOOP_for_if_2_for_for_if_aelse_acc_nl[8:0];
  assign LOAD_LOOP_for_if_2_for_for_if_aelse_acc_itm_8 = readslicef_9_1_8(LOAD_LOOP_for_if_2_for_for_if_aelse_acc_nl);
  assign nl_operator_8_false_6_acc_nl = conv_u2s_4_5(LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1[4:1])
      + 5'b10111;
  assign operator_8_false_6_acc_nl = nl_operator_8_false_6_acc_nl[4:0];
  assign operator_8_false_6_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_6_acc_nl);
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d = LOAD_LOOP_for_if_2_for_for_if_mux_rmff;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d = LOAD_LOOP_for_if_2_for_for_else_index_in_mux_rmff;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d = LOAD_LOOP_for_if_2_for_for_if_index_in_mux_rmff;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff = LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_iff;
  assign LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d =
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign or_dcpl_395 = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 | LOAD_LOOP_for_if_2_for_nor_tmp_1
      | LOAD_LOOP_for_if_2_for_and_199_cse;
  assign or_dcpl_401 = LOAD_LOOP_for_if_2_for_nor_tmp_1 | LOAD_LOOP_for_if_2_for_or_tmp_1
      | LOAD_LOOP_for_if_2_for_and_180_cse_1;
  assign nor_794_nl = ~(nor_178_cse | LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign or_2906_nl = (~ LOAD_BATCH_LOOP_stage_v_1) | LOAD_BATCH_LOOP_asn_itm_1;
  assign mux_tmp = MUX_s_1_2_2(nor_794_nl, exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2,
      or_2906_nl);
  assign and_3316_cse = (mux_tmp | LOAD_LOOP_for_LOAD_LOOP_nand_cse) & (fsm_output[2]);
  assign and_3318_cse = (~ mux_tmp) & and_3266_cse & (fsm_output[2]);
  assign and_3338_cse = (conf_info_crt_sva_231_0[98]) & (fsm_output[2]);
  assign or_tmp_2431 = (conf_info_crt_sva_231_0[97]) & (fsm_output[2]);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_idat_15_0 <= 16'b0000000000000000;
    end
    else if ( core_wen & (or_tmp_1480 | or_tmp_1481 | dma_read_ctrl_rsci_idat_15_0_mx0c2)
        ) begin
      dma_read_ctrl_rsci_idat_15_0 <= MUX1HOT_v_16_3_2((z_out_10[15:0]), LOAD_LOOP_for_ac_int_cctor_lpi_2,
          LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2, {LOAD_CTRL_LOOP1_or_nl , LOAD_CTRL_LOOP1_and_2_nl
          , dma_read_ctrl_rsci_idat_15_0_mx0c2});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( core_wen & (or_tmp_1480 | dma_read_ctrl_rsci_idat_47_32_mx0c1) ) begin
      dma_read_ctrl_rsci_idat_47_32 <= MUX_v_16_2_2(batch_size_mul_4_cse_sva, batch_size_mul_1_cse_sva,
          dma_read_ctrl_rsci_idat_47_32_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_36 & (fsm_output[2])) | plm_kernel_rsci_idat_31_0_mx0c1)
        ) begin
      plm_kernel_rsci_idat_31_0 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt, LOAD_BATCH_LOOP_plm_tmp_f_data_0_sva,
          plm_kernel_rsci_idat_31_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_47 & (fsm_output[2])) | plm_kernel_rsci_idat_63_32_mx0c1)
        ) begin
      plm_kernel_rsci_idat_63_32 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt, LOAD_BATCH_LOOP_plm_tmp_f_data_1_sva,
          plm_kernel_rsci_idat_63_32_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_51 & (fsm_output[2])) | plm_kernel_rsci_idat_95_64_mx0c1)
        ) begin
      plm_kernel_rsci_idat_95_64 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt, LOAD_BATCH_LOOP_plm_tmp_f_data_2_sva,
          plm_kernel_rsci_idat_95_64_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_127_96 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_54 & (fsm_output[2])) | plm_kernel_rsci_idat_127_96_mx0c1)
        ) begin
      plm_kernel_rsci_idat_127_96 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt, LOAD_BATCH_LOOP_plm_tmp_f_data_3_sva,
          plm_kernel_rsci_idat_127_96_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_159_128 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_58 & (fsm_output[2])) | plm_kernel_rsci_idat_159_128_mx0c1)
        ) begin
      plm_kernel_rsci_idat_159_128 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_4_sva, plm_kernel_rsci_idat_159_128_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_191_160 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_62 & (fsm_output[2])) | plm_kernel_rsci_idat_191_160_mx0c1)
        ) begin
      plm_kernel_rsci_idat_191_160 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_5_sva, plm_kernel_rsci_idat_191_160_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_223_192 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_65 & (fsm_output[2])) | plm_kernel_rsci_idat_223_192_mx0c1)
        ) begin
      plm_kernel_rsci_idat_223_192 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_6_sva, plm_kernel_rsci_idat_223_192_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_255_224 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_41 & and_dcpl_68 & (fsm_output[2])) | plm_kernel_rsci_idat_255_224_mx0c1)
        ) begin
      plm_kernel_rsci_idat_255_224 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_7_sva, plm_kernel_rsci_idat_255_224_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_287_256 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_36 & (fsm_output[2])) | plm_kernel_rsci_idat_287_256_mx0c1)
        ) begin
      plm_kernel_rsci_idat_287_256 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_8_sva, plm_kernel_rsci_idat_287_256_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_319_288 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_47 & (fsm_output[2])) | plm_kernel_rsci_idat_319_288_mx0c1)
        ) begin
      plm_kernel_rsci_idat_319_288 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_9_sva, plm_kernel_rsci_idat_319_288_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_351_320 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_51 & (fsm_output[2])) | plm_kernel_rsci_idat_351_320_mx0c1)
        ) begin
      plm_kernel_rsci_idat_351_320 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_10_sva, plm_kernel_rsci_idat_351_320_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_383_352 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_54 & (fsm_output[2])) | plm_kernel_rsci_idat_383_352_mx0c1)
        ) begin
      plm_kernel_rsci_idat_383_352 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_11_sva, plm_kernel_rsci_idat_383_352_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_415_384 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_58 & (fsm_output[2])) | plm_kernel_rsci_idat_415_384_mx0c1)
        ) begin
      plm_kernel_rsci_idat_415_384 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_12_sva, plm_kernel_rsci_idat_415_384_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_447_416 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_62 & (fsm_output[2])) | plm_kernel_rsci_idat_447_416_mx0c1)
        ) begin
      plm_kernel_rsci_idat_447_416 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_13_sva, plm_kernel_rsci_idat_447_416_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_479_448 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_65 & (fsm_output[2])) | plm_kernel_rsci_idat_479_448_mx0c1)
        ) begin
      plm_kernel_rsci_idat_479_448 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_14_sva, plm_kernel_rsci_idat_479_448_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_511_480 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_72 & and_dcpl_68 & (fsm_output[2])) | plm_kernel_rsci_idat_511_480_mx0c1)
        ) begin
      plm_kernel_rsci_idat_511_480 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_15_sva, plm_kernel_rsci_idat_511_480_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_543_512 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_36 & (fsm_output[2])) | plm_kernel_rsci_idat_543_512_mx0c1)
        ) begin
      plm_kernel_rsci_idat_543_512 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_16_sva, plm_kernel_rsci_idat_543_512_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_575_544 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_47 & (fsm_output[2])) | plm_kernel_rsci_idat_575_544_mx0c1)
        ) begin
      plm_kernel_rsci_idat_575_544 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_17_sva, plm_kernel_rsci_idat_575_544_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_607_576 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_51 & (fsm_output[2])) | plm_kernel_rsci_idat_607_576_mx0c1)
        ) begin
      plm_kernel_rsci_idat_607_576 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_18_sva, plm_kernel_rsci_idat_607_576_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_639_608 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_54 & (fsm_output[2])) | plm_kernel_rsci_idat_639_608_mx0c1)
        ) begin
      plm_kernel_rsci_idat_639_608 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_19_sva, plm_kernel_rsci_idat_639_608_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_671_640 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_58 & (fsm_output[2])) | plm_kernel_rsci_idat_671_640_mx0c1)
        ) begin
      plm_kernel_rsci_idat_671_640 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_20_sva, plm_kernel_rsci_idat_671_640_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_703_672 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_62 & (fsm_output[2])) | plm_kernel_rsci_idat_703_672_mx0c1)
        ) begin
      plm_kernel_rsci_idat_703_672 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_21_sva, plm_kernel_rsci_idat_703_672_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_735_704 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_65 & (fsm_output[2])) | plm_kernel_rsci_idat_735_704_mx0c1)
        ) begin
      plm_kernel_rsci_idat_735_704 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_22_sva, plm_kernel_rsci_idat_735_704_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_767_736 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_91 & and_dcpl_68 & (fsm_output[2])) | plm_kernel_rsci_idat_767_736_mx0c1)
        ) begin
      plm_kernel_rsci_idat_767_736 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_23_sva, plm_kernel_rsci_idat_767_736_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_799_768 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_36 & (fsm_output[2])) | plm_kernel_rsci_idat_799_768_mx0c1)
        ) begin
      plm_kernel_rsci_idat_799_768 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_24_sva, plm_kernel_rsci_idat_799_768_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_831_800 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_47 & (fsm_output[2])) | plm_kernel_rsci_idat_831_800_mx0c1)
        ) begin
      plm_kernel_rsci_idat_831_800 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_25_sva, plm_kernel_rsci_idat_831_800_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_863_832 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_51 & (fsm_output[2])) | plm_kernel_rsci_idat_863_832_mx0c1)
        ) begin
      plm_kernel_rsci_idat_863_832 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_26_sva, plm_kernel_rsci_idat_863_832_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_895_864 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_54 & (fsm_output[2])) | plm_kernel_rsci_idat_895_864_mx0c1)
        ) begin
      plm_kernel_rsci_idat_895_864 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_27_sva, plm_kernel_rsci_idat_895_864_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_927_896 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_58 & (fsm_output[2])) | plm_kernel_rsci_idat_927_896_mx0c1)
        ) begin
      plm_kernel_rsci_idat_927_896 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_28_sva, plm_kernel_rsci_idat_927_896_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_959_928 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_62 & (fsm_output[2])) | plm_kernel_rsci_idat_959_928_mx0c1)
        ) begin
      plm_kernel_rsci_idat_959_928 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_29_sva, plm_kernel_rsci_idat_959_928_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_991_960 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_65 & (fsm_output[2])) | plm_kernel_rsci_idat_991_960_mx0c1)
        ) begin
      plm_kernel_rsci_idat_991_960 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_30_sva, plm_kernel_rsci_idat_991_960_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1023_992 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_108 & and_dcpl_68 & (fsm_output[2])) | plm_kernel_rsci_idat_1023_992_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1023_992 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_31_sva, plm_kernel_rsci_idat_1023_992_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1055_1024 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_36 & (fsm_output[2])) | plm_kernel_rsci_idat_1055_1024_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1055_1024 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_32_sva, plm_kernel_rsci_idat_1055_1024_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1087_1056 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_47 & (fsm_output[2])) | plm_kernel_rsci_idat_1087_1056_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1087_1056 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_33_sva, plm_kernel_rsci_idat_1087_1056_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1119_1088 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_51 & (fsm_output[2])) | plm_kernel_rsci_idat_1119_1088_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1119_1088 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_34_sva, plm_kernel_rsci_idat_1119_1088_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1151_1120 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_54 & (fsm_output[2])) | plm_kernel_rsci_idat_1151_1120_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1151_1120 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_35_sva, plm_kernel_rsci_idat_1151_1120_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1183_1152 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_58 & (fsm_output[2])) | plm_kernel_rsci_idat_1183_1152_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1183_1152 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_36_sva, plm_kernel_rsci_idat_1183_1152_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1215_1184 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_62 & (fsm_output[2])) | plm_kernel_rsci_idat_1215_1184_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1215_1184 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_37_sva, plm_kernel_rsci_idat_1215_1184_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1247_1216 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_65 & (fsm_output[2])) | plm_kernel_rsci_idat_1247_1216_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1247_1216 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_38_sva, plm_kernel_rsci_idat_1247_1216_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1279_1248 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_127 & and_dcpl_68 & (fsm_output[2])) | plm_kernel_rsci_idat_1279_1248_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1279_1248 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_39_sva, plm_kernel_rsci_idat_1279_1248_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1311_1280 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_36 & (fsm_output[2])) | plm_kernel_rsci_idat_1311_1280_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1311_1280 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_40_sva, plm_kernel_rsci_idat_1311_1280_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1343_1312 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_47 & (fsm_output[2])) | plm_kernel_rsci_idat_1343_1312_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1343_1312 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_41_sva, plm_kernel_rsci_idat_1343_1312_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1375_1344 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_51 & (fsm_output[2])) | plm_kernel_rsci_idat_1375_1344_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1375_1344 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_42_sva, plm_kernel_rsci_idat_1375_1344_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1407_1376 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_54 & (fsm_output[2])) | plm_kernel_rsci_idat_1407_1376_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1407_1376 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_43_sva, plm_kernel_rsci_idat_1407_1376_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1439_1408 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_58 & (fsm_output[2])) | plm_kernel_rsci_idat_1439_1408_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1439_1408 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_44_sva, plm_kernel_rsci_idat_1439_1408_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1471_1440 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_62 & (fsm_output[2])) | plm_kernel_rsci_idat_1471_1440_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1471_1440 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_45_sva, plm_kernel_rsci_idat_1471_1440_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1503_1472 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_65 & (fsm_output[2])) | plm_kernel_rsci_idat_1503_1472_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1503_1472 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_46_sva, plm_kernel_rsci_idat_1503_1472_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1535_1504 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_144 & and_dcpl_68 & (fsm_output[2])) | plm_kernel_rsci_idat_1535_1504_mx0c1)
        ) begin
      plm_kernel_rsci_idat_1535_1504 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_47_sva, plm_kernel_rsci_idat_1535_1504_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_kernel_rsci_idat_1567_1536 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_40 & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b11)
        & (~ (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0])) & and_dcpl_36
        & (fsm_output[2])) | plm_kernel_rsci_idat_1567_1536_mx0c1) ) begin
      plm_kernel_rsci_idat_1567_1536 <= MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
          LOAD_BATCH_LOOP_plm_tmp_f_data_48_sva, plm_kernel_rsci_idat_1567_1536_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_169 & (fsm_output[2]))
        | buf_linear_rsci_idat_31_0_mx0c1) ) begin
      buf_linear_rsci_idat_31_0 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_0_sva, buf_linear_rsci_idat_31_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_169 & (fsm_output[2]))
        | buf_linear_rsci_idat_63_32_mx0c1) ) begin
      buf_linear_rsci_idat_63_32 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_1_sva, buf_linear_rsci_idat_63_32_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_95_64 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_169 & (fsm_output[2]))
        | buf_linear_rsci_idat_95_64_mx0c1) ) begin
      buf_linear_rsci_idat_95_64 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_2_sva, buf_linear_rsci_idat_95_64_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_127_96 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_169 & (fsm_output[2]))
        | buf_linear_rsci_idat_127_96_mx0c1) ) begin
      buf_linear_rsci_idat_127_96 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_3_sva, buf_linear_rsci_idat_127_96_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_159_128 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_206 & (fsm_output[2]))
        | buf_linear_rsci_idat_159_128_mx0c1) ) begin
      buf_linear_rsci_idat_159_128 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_4_sva, buf_linear_rsci_idat_159_128_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_191_160 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_206 & (fsm_output[2]))
        | buf_linear_rsci_idat_191_160_mx0c1) ) begin
      buf_linear_rsci_idat_191_160 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_5_sva, buf_linear_rsci_idat_191_160_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_223_192 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_206 & (fsm_output[2]))
        | buf_linear_rsci_idat_223_192_mx0c1) ) begin
      buf_linear_rsci_idat_223_192 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_6_sva, buf_linear_rsci_idat_223_192_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_255_224 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_206 & (fsm_output[2]))
        | buf_linear_rsci_idat_255_224_mx0c1) ) begin
      buf_linear_rsci_idat_255_224 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_7_sva, buf_linear_rsci_idat_255_224_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_287_256 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_224 & (fsm_output[2]))
        | buf_linear_rsci_idat_287_256_mx0c1) ) begin
      buf_linear_rsci_idat_287_256 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_8_sva, buf_linear_rsci_idat_287_256_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_319_288 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_224 & (fsm_output[2]))
        | buf_linear_rsci_idat_319_288_mx0c1) ) begin
      buf_linear_rsci_idat_319_288 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_9_sva, buf_linear_rsci_idat_319_288_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_351_320 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_224 & (fsm_output[2]))
        | buf_linear_rsci_idat_351_320_mx0c1) ) begin
      buf_linear_rsci_idat_351_320 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_10_sva, buf_linear_rsci_idat_351_320_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_383_352 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_224 & (fsm_output[2]))
        | buf_linear_rsci_idat_383_352_mx0c1) ) begin
      buf_linear_rsci_idat_383_352 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_11_sva, buf_linear_rsci_idat_383_352_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_415_384 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_242 & (fsm_output[2]))
        | buf_linear_rsci_idat_415_384_mx0c1) ) begin
      buf_linear_rsci_idat_415_384 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_12_sva, buf_linear_rsci_idat_415_384_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_447_416 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_242 & (fsm_output[2]))
        | buf_linear_rsci_idat_447_416_mx0c1) ) begin
      buf_linear_rsci_idat_447_416 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_13_sva, buf_linear_rsci_idat_447_416_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_479_448 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_242 & (fsm_output[2]))
        | buf_linear_rsci_idat_479_448_mx0c1) ) begin
      buf_linear_rsci_idat_479_448 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_14_sva, buf_linear_rsci_idat_479_448_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_511_480 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_242 & (fsm_output[2]))
        | buf_linear_rsci_idat_511_480_mx0c1) ) begin
      buf_linear_rsci_idat_511_480 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_15_sva, buf_linear_rsci_idat_511_480_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_543_512 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_260 & (fsm_output[2]))
        | buf_linear_rsci_idat_543_512_mx0c1) ) begin
      buf_linear_rsci_idat_543_512 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_16_sva, buf_linear_rsci_idat_543_512_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_575_544 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_260 & (fsm_output[2]))
        | buf_linear_rsci_idat_575_544_mx0c1) ) begin
      buf_linear_rsci_idat_575_544 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_0_17_sva, buf_linear_rsci_idat_575_544_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_607_576 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_260 & (fsm_output[2]))
        | buf_linear_rsci_idat_607_576_mx0c1) ) begin
      buf_linear_rsci_idat_607_576 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_0_sva, buf_linear_rsci_idat_607_576_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_639_608 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_260 & (fsm_output[2]))
        | buf_linear_rsci_idat_639_608_mx0c1) ) begin
      buf_linear_rsci_idat_639_608 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_1_sva, buf_linear_rsci_idat_639_608_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_671_640 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_277 & (fsm_output[2]))
        | buf_linear_rsci_idat_671_640_mx0c1) ) begin
      buf_linear_rsci_idat_671_640 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_2_sva, buf_linear_rsci_idat_671_640_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_703_672 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_277 & (fsm_output[2]))
        | buf_linear_rsci_idat_703_672_mx0c1) ) begin
      buf_linear_rsci_idat_703_672 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_3_sva, buf_linear_rsci_idat_703_672_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_735_704 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_277 & (fsm_output[2]))
        | buf_linear_rsci_idat_735_704_mx0c1) ) begin
      buf_linear_rsci_idat_735_704 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_4_sva, buf_linear_rsci_idat_735_704_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_767_736 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_277 & (fsm_output[2]))
        | buf_linear_rsci_idat_767_736_mx0c1) ) begin
      buf_linear_rsci_idat_767_736 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_5_sva, buf_linear_rsci_idat_767_736_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_799_768 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_294 & (fsm_output[2]))
        | buf_linear_rsci_idat_799_768_mx0c1) ) begin
      buf_linear_rsci_idat_799_768 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_6_sva, buf_linear_rsci_idat_799_768_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_831_800 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_294 & (fsm_output[2]))
        | buf_linear_rsci_idat_831_800_mx0c1) ) begin
      buf_linear_rsci_idat_831_800 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_7_sva, buf_linear_rsci_idat_831_800_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_863_832 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_294 & (fsm_output[2]))
        | buf_linear_rsci_idat_863_832_mx0c1) ) begin
      buf_linear_rsci_idat_863_832 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_8_sva, buf_linear_rsci_idat_863_832_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_895_864 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_294 & (fsm_output[2]))
        | buf_linear_rsci_idat_895_864_mx0c1) ) begin
      buf_linear_rsci_idat_895_864 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_9_sva, buf_linear_rsci_idat_895_864_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_927_896 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_311 & (fsm_output[2]))
        | buf_linear_rsci_idat_927_896_mx0c1) ) begin
      buf_linear_rsci_idat_927_896 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_10_sva, buf_linear_rsci_idat_927_896_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_959_928 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_311 & (fsm_output[2]))
        | buf_linear_rsci_idat_959_928_mx0c1) ) begin
      buf_linear_rsci_idat_959_928 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_11_sva, buf_linear_rsci_idat_959_928_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_991_960 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_311 & (fsm_output[2]))
        | buf_linear_rsci_idat_991_960_mx0c1) ) begin
      buf_linear_rsci_idat_991_960 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_12_sva, buf_linear_rsci_idat_991_960_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1023_992 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_311 & (fsm_output[2]))
        | buf_linear_rsci_idat_1023_992_mx0c1) ) begin
      buf_linear_rsci_idat_1023_992 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_13_sva, buf_linear_rsci_idat_1023_992_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1055_1024 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_330 & (fsm_output[2]))
        | buf_linear_rsci_idat_1055_1024_mx0c1) ) begin
      buf_linear_rsci_idat_1055_1024 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_14_sva, buf_linear_rsci_idat_1055_1024_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1087_1056 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_330 & (fsm_output[2]))
        | buf_linear_rsci_idat_1087_1056_mx0c1) ) begin
      buf_linear_rsci_idat_1087_1056 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_15_sva, buf_linear_rsci_idat_1087_1056_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1119_1088 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_330 & (fsm_output[2]))
        | buf_linear_rsci_idat_1119_1088_mx0c1) ) begin
      buf_linear_rsci_idat_1119_1088 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_16_sva, buf_linear_rsci_idat_1119_1088_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1151_1120 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_330 & (fsm_output[2]))
        | buf_linear_rsci_idat_1151_1120_mx0c1) ) begin
      buf_linear_rsci_idat_1151_1120 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_1_17_sva, buf_linear_rsci_idat_1151_1120_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1183_1152 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_347 & (fsm_output[2]))
        | buf_linear_rsci_idat_1183_1152_mx0c1) ) begin
      buf_linear_rsci_idat_1183_1152 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_0_sva, buf_linear_rsci_idat_1183_1152_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1215_1184 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_347 & (fsm_output[2]))
        | buf_linear_rsci_idat_1215_1184_mx0c1) ) begin
      buf_linear_rsci_idat_1215_1184 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_1_sva, buf_linear_rsci_idat_1215_1184_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1247_1216 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_347 & (fsm_output[2]))
        | buf_linear_rsci_idat_1247_1216_mx0c1) ) begin
      buf_linear_rsci_idat_1247_1216 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_2_sva, buf_linear_rsci_idat_1247_1216_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1279_1248 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_347 & (fsm_output[2]))
        | buf_linear_rsci_idat_1279_1248_mx0c1) ) begin
      buf_linear_rsci_idat_1279_1248 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_3_sva, buf_linear_rsci_idat_1279_1248_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1311_1280 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_364 & (fsm_output[2]))
        | buf_linear_rsci_idat_1311_1280_mx0c1) ) begin
      buf_linear_rsci_idat_1311_1280 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_4_sva, buf_linear_rsci_idat_1311_1280_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1343_1312 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_364 & (fsm_output[2]))
        | buf_linear_rsci_idat_1343_1312_mx0c1) ) begin
      buf_linear_rsci_idat_1343_1312 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_5_sva, buf_linear_rsci_idat_1343_1312_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1375_1344 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_364 & (fsm_output[2]))
        | buf_linear_rsci_idat_1375_1344_mx0c1) ) begin
      buf_linear_rsci_idat_1375_1344 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_6_sva, buf_linear_rsci_idat_1375_1344_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1407_1376 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_364 & (fsm_output[2]))
        | buf_linear_rsci_idat_1407_1376_mx0c1) ) begin
      buf_linear_rsci_idat_1407_1376 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_7_sva, buf_linear_rsci_idat_1407_1376_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1439_1408 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_381 & (fsm_output[2]))
        | buf_linear_rsci_idat_1439_1408_mx0c1) ) begin
      buf_linear_rsci_idat_1439_1408 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_8_sva, buf_linear_rsci_idat_1439_1408_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1471_1440 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_381 & (fsm_output[2]))
        | buf_linear_rsci_idat_1471_1440_mx0c1) ) begin
      buf_linear_rsci_idat_1471_1440 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_9_sva, buf_linear_rsci_idat_1471_1440_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1503_1472 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_381 & (fsm_output[2]))
        | buf_linear_rsci_idat_1503_1472_mx0c1) ) begin
      buf_linear_rsci_idat_1503_1472 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_10_sva, buf_linear_rsci_idat_1503_1472_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1535_1504 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_381 & (fsm_output[2]))
        | buf_linear_rsci_idat_1535_1504_mx0c1) ) begin
      buf_linear_rsci_idat_1535_1504 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_11_sva, buf_linear_rsci_idat_1535_1504_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1567_1536 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_399 & (fsm_output[2]))
        | buf_linear_rsci_idat_1567_1536_mx0c1) ) begin
      buf_linear_rsci_idat_1567_1536 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_12_sva, buf_linear_rsci_idat_1567_1536_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1599_1568 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_399 & (fsm_output[2]))
        | buf_linear_rsci_idat_1599_1568_mx0c1) ) begin
      buf_linear_rsci_idat_1599_1568 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_13_sva, buf_linear_rsci_idat_1599_1568_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1631_1600 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_399 & (fsm_output[2]))
        | buf_linear_rsci_idat_1631_1600_mx0c1) ) begin
      buf_linear_rsci_idat_1631_1600 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_14_sva, buf_linear_rsci_idat_1631_1600_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1663_1632 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_399 & (fsm_output[2]))
        | buf_linear_rsci_idat_1663_1632_mx0c1) ) begin
      buf_linear_rsci_idat_1663_1632 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_15_sva, buf_linear_rsci_idat_1663_1632_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1695_1664 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_416 & (fsm_output[2]))
        | buf_linear_rsci_idat_1695_1664_mx0c1) ) begin
      buf_linear_rsci_idat_1695_1664 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_16_sva, buf_linear_rsci_idat_1695_1664_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1727_1696 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_416 & (fsm_output[2]))
        | buf_linear_rsci_idat_1727_1696_mx0c1) ) begin
      buf_linear_rsci_idat_1727_1696 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_2_17_sva, buf_linear_rsci_idat_1727_1696_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1759_1728 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_416 & (fsm_output[2]))
        | buf_linear_rsci_idat_1759_1728_mx0c1) ) begin
      buf_linear_rsci_idat_1759_1728 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_0_sva, buf_linear_rsci_idat_1759_1728_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1791_1760 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_416 & (fsm_output[2]))
        | buf_linear_rsci_idat_1791_1760_mx0c1) ) begin
      buf_linear_rsci_idat_1791_1760 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_1_sva, buf_linear_rsci_idat_1791_1760_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1823_1792 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_433 & (fsm_output[2]))
        | buf_linear_rsci_idat_1823_1792_mx0c1) ) begin
      buf_linear_rsci_idat_1823_1792 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_2_sva, buf_linear_rsci_idat_1823_1792_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1855_1824 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_433 & (fsm_output[2]))
        | buf_linear_rsci_idat_1855_1824_mx0c1) ) begin
      buf_linear_rsci_idat_1855_1824 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_3_sva, buf_linear_rsci_idat_1855_1824_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1887_1856 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_433 & (fsm_output[2]))
        | buf_linear_rsci_idat_1887_1856_mx0c1) ) begin
      buf_linear_rsci_idat_1887_1856 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_4_sva, buf_linear_rsci_idat_1887_1856_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1919_1888 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_433 & (fsm_output[2]))
        | buf_linear_rsci_idat_1919_1888_mx0c1) ) begin
      buf_linear_rsci_idat_1919_1888 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_5_sva, buf_linear_rsci_idat_1919_1888_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1951_1920 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_450 & (fsm_output[2]))
        | buf_linear_rsci_idat_1951_1920_mx0c1) ) begin
      buf_linear_rsci_idat_1951_1920 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_6_sva, buf_linear_rsci_idat_1951_1920_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_1983_1952 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_450 & (fsm_output[2]))
        | buf_linear_rsci_idat_1983_1952_mx0c1) ) begin
      buf_linear_rsci_idat_1983_1952 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_7_sva, buf_linear_rsci_idat_1983_1952_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2015_1984 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_450 & (fsm_output[2]))
        | buf_linear_rsci_idat_2015_1984_mx0c1) ) begin
      buf_linear_rsci_idat_2015_1984 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_8_sva, buf_linear_rsci_idat_2015_1984_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2047_2016 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_450 & (fsm_output[2]))
        | buf_linear_rsci_idat_2047_2016_mx0c1) ) begin
      buf_linear_rsci_idat_2047_2016 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_9_sva, buf_linear_rsci_idat_2047_2016_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2079_2048 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_469 & (fsm_output[2]))
        | buf_linear_rsci_idat_2079_2048_mx0c1) ) begin
      buf_linear_rsci_idat_2079_2048 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_10_sva, buf_linear_rsci_idat_2079_2048_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2111_2080 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_469 & (fsm_output[2]))
        | buf_linear_rsci_idat_2111_2080_mx0c1) ) begin
      buf_linear_rsci_idat_2111_2080 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_11_sva, buf_linear_rsci_idat_2111_2080_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2143_2112 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_469 & (fsm_output[2]))
        | buf_linear_rsci_idat_2143_2112_mx0c1) ) begin
      buf_linear_rsci_idat_2143_2112 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_12_sva, buf_linear_rsci_idat_2143_2112_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2175_2144 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_469 & (fsm_output[2]))
        | buf_linear_rsci_idat_2175_2144_mx0c1) ) begin
      buf_linear_rsci_idat_2175_2144 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_13_sva, buf_linear_rsci_idat_2175_2144_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2207_2176 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_486 & (fsm_output[2]))
        | buf_linear_rsci_idat_2207_2176_mx0c1) ) begin
      buf_linear_rsci_idat_2207_2176 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_14_sva, buf_linear_rsci_idat_2207_2176_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2239_2208 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_486 & (fsm_output[2]))
        | buf_linear_rsci_idat_2239_2208_mx0c1) ) begin
      buf_linear_rsci_idat_2239_2208 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_15_sva, buf_linear_rsci_idat_2239_2208_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2271_2240 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_486 & (fsm_output[2]))
        | buf_linear_rsci_idat_2271_2240_mx0c1) ) begin
      buf_linear_rsci_idat_2271_2240 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_16_sva, buf_linear_rsci_idat_2271_2240_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2303_2272 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_486 & (fsm_output[2]))
        | buf_linear_rsci_idat_2303_2272_mx0c1) ) begin
      buf_linear_rsci_idat_2303_2272 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_3_17_sva, buf_linear_rsci_idat_2303_2272_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2335_2304 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_503 & (fsm_output[2]))
        | buf_linear_rsci_idat_2335_2304_mx0c1) ) begin
      buf_linear_rsci_idat_2335_2304 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_0_sva, buf_linear_rsci_idat_2335_2304_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2367_2336 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_503 & (fsm_output[2]))
        | buf_linear_rsci_idat_2367_2336_mx0c1) ) begin
      buf_linear_rsci_idat_2367_2336 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_1_sva, buf_linear_rsci_idat_2367_2336_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2399_2368 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_503 & (fsm_output[2]))
        | buf_linear_rsci_idat_2399_2368_mx0c1) ) begin
      buf_linear_rsci_idat_2399_2368 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_2_sva, buf_linear_rsci_idat_2399_2368_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2431_2400 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_503 & (fsm_output[2]))
        | buf_linear_rsci_idat_2431_2400_mx0c1) ) begin
      buf_linear_rsci_idat_2431_2400 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_3_sva, buf_linear_rsci_idat_2431_2400_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2463_2432 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_520 & (fsm_output[2]))
        | buf_linear_rsci_idat_2463_2432_mx0c1) ) begin
      buf_linear_rsci_idat_2463_2432 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_4_sva, buf_linear_rsci_idat_2463_2432_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2495_2464 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_520 & (fsm_output[2]))
        | buf_linear_rsci_idat_2495_2464_mx0c1) ) begin
      buf_linear_rsci_idat_2495_2464 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_5_sva, buf_linear_rsci_idat_2495_2464_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2527_2496 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_520 & (fsm_output[2]))
        | buf_linear_rsci_idat_2527_2496_mx0c1) ) begin
      buf_linear_rsci_idat_2527_2496 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_6_sva, buf_linear_rsci_idat_2527_2496_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2559_2528 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_520 & (fsm_output[2]))
        | buf_linear_rsci_idat_2559_2528_mx0c1) ) begin
      buf_linear_rsci_idat_2559_2528 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_7_sva, buf_linear_rsci_idat_2559_2528_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2591_2560 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_538 & (fsm_output[2]))
        | buf_linear_rsci_idat_2591_2560_mx0c1) ) begin
      buf_linear_rsci_idat_2591_2560 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_8_sva, buf_linear_rsci_idat_2591_2560_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2623_2592 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_538 & (fsm_output[2]))
        | buf_linear_rsci_idat_2623_2592_mx0c1) ) begin
      buf_linear_rsci_idat_2623_2592 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_9_sva, buf_linear_rsci_idat_2623_2592_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2655_2624 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_538 & (fsm_output[2]))
        | buf_linear_rsci_idat_2655_2624_mx0c1) ) begin
      buf_linear_rsci_idat_2655_2624 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_10_sva, buf_linear_rsci_idat_2655_2624_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2687_2656 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_538 & (fsm_output[2]))
        | buf_linear_rsci_idat_2687_2656_mx0c1) ) begin
      buf_linear_rsci_idat_2687_2656 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_11_sva, buf_linear_rsci_idat_2687_2656_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2719_2688 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_555 & (fsm_output[2]))
        | buf_linear_rsci_idat_2719_2688_mx0c1) ) begin
      buf_linear_rsci_idat_2719_2688 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_12_sva, buf_linear_rsci_idat_2719_2688_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2751_2720 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_555 & (fsm_output[2]))
        | buf_linear_rsci_idat_2751_2720_mx0c1) ) begin
      buf_linear_rsci_idat_2751_2720 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_13_sva, buf_linear_rsci_idat_2751_2720_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2783_2752 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_555 & (fsm_output[2]))
        | buf_linear_rsci_idat_2783_2752_mx0c1) ) begin
      buf_linear_rsci_idat_2783_2752 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_14_sva, buf_linear_rsci_idat_2783_2752_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2815_2784 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_555 & (fsm_output[2]))
        | buf_linear_rsci_idat_2815_2784_mx0c1) ) begin
      buf_linear_rsci_idat_2815_2784 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_15_sva, buf_linear_rsci_idat_2815_2784_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2847_2816 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_572 & (fsm_output[2]))
        | buf_linear_rsci_idat_2847_2816_mx0c1) ) begin
      buf_linear_rsci_idat_2847_2816 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_16_sva, buf_linear_rsci_idat_2847_2816_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2879_2848 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_572 & (fsm_output[2]))
        | buf_linear_rsci_idat_2879_2848_mx0c1) ) begin
      buf_linear_rsci_idat_2879_2848 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_4_17_sva, buf_linear_rsci_idat_2879_2848_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2911_2880 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_572 & (fsm_output[2]))
        | buf_linear_rsci_idat_2911_2880_mx0c1) ) begin
      buf_linear_rsci_idat_2911_2880 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_0_sva, buf_linear_rsci_idat_2911_2880_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2943_2912 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_572 & (fsm_output[2]))
        | buf_linear_rsci_idat_2943_2912_mx0c1) ) begin
      buf_linear_rsci_idat_2943_2912 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_1_sva, buf_linear_rsci_idat_2943_2912_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_2975_2944 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_589 & (fsm_output[2]))
        | buf_linear_rsci_idat_2975_2944_mx0c1) ) begin
      buf_linear_rsci_idat_2975_2944 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_2_sva, buf_linear_rsci_idat_2975_2944_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3007_2976 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_589 & (fsm_output[2]))
        | buf_linear_rsci_idat_3007_2976_mx0c1) ) begin
      buf_linear_rsci_idat_3007_2976 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_3_sva, buf_linear_rsci_idat_3007_2976_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3039_3008 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_589 & (fsm_output[2]))
        | buf_linear_rsci_idat_3039_3008_mx0c1) ) begin
      buf_linear_rsci_idat_3039_3008 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_4_sva, buf_linear_rsci_idat_3039_3008_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3071_3040 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_589 & (fsm_output[2]))
        | buf_linear_rsci_idat_3071_3040_mx0c1) ) begin
      buf_linear_rsci_idat_3071_3040 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_5_sva, buf_linear_rsci_idat_3071_3040_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3103_3072 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_608 & (fsm_output[2]))
        | buf_linear_rsci_idat_3103_3072_mx0c1) ) begin
      buf_linear_rsci_idat_3103_3072 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_6_sva, buf_linear_rsci_idat_3103_3072_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3135_3104 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_608 & (fsm_output[2]))
        | buf_linear_rsci_idat_3135_3104_mx0c1) ) begin
      buf_linear_rsci_idat_3135_3104 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_7_sva, buf_linear_rsci_idat_3135_3104_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3167_3136 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_608 & (fsm_output[2]))
        | buf_linear_rsci_idat_3167_3136_mx0c1) ) begin
      buf_linear_rsci_idat_3167_3136 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_8_sva, buf_linear_rsci_idat_3167_3136_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3199_3168 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_608 & (fsm_output[2]))
        | buf_linear_rsci_idat_3199_3168_mx0c1) ) begin
      buf_linear_rsci_idat_3199_3168 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_9_sva, buf_linear_rsci_idat_3199_3168_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3231_3200 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_625 & (fsm_output[2]))
        | buf_linear_rsci_idat_3231_3200_mx0c1) ) begin
      buf_linear_rsci_idat_3231_3200 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_10_sva, buf_linear_rsci_idat_3231_3200_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3263_3232 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_625 & (fsm_output[2]))
        | buf_linear_rsci_idat_3263_3232_mx0c1) ) begin
      buf_linear_rsci_idat_3263_3232 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_11_sva, buf_linear_rsci_idat_3263_3232_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3295_3264 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_625 & (fsm_output[2]))
        | buf_linear_rsci_idat_3295_3264_mx0c1) ) begin
      buf_linear_rsci_idat_3295_3264 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_12_sva, buf_linear_rsci_idat_3295_3264_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3327_3296 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_625 & (fsm_output[2]))
        | buf_linear_rsci_idat_3327_3296_mx0c1) ) begin
      buf_linear_rsci_idat_3327_3296 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_13_sva, buf_linear_rsci_idat_3327_3296_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3359_3328 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_642 & (fsm_output[2]))
        | buf_linear_rsci_idat_3359_3328_mx0c1) ) begin
      buf_linear_rsci_idat_3359_3328 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_14_sva, buf_linear_rsci_idat_3359_3328_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3391_3360 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_642 & (fsm_output[2]))
        | buf_linear_rsci_idat_3391_3360_mx0c1) ) begin
      buf_linear_rsci_idat_3391_3360 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_15_sva, buf_linear_rsci_idat_3391_3360_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3423_3392 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_642 & (fsm_output[2]))
        | buf_linear_rsci_idat_3423_3392_mx0c1) ) begin
      buf_linear_rsci_idat_3423_3392 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_16_sva, buf_linear_rsci_idat_3423_3392_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3455_3424 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_642 & (fsm_output[2]))
        | buf_linear_rsci_idat_3455_3424_mx0c1) ) begin
      buf_linear_rsci_idat_3455_3424 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_5_17_sva, buf_linear_rsci_idat_3455_3424_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3487_3456 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_659 & (fsm_output[2]))
        | buf_linear_rsci_idat_3487_3456_mx0c1) ) begin
      buf_linear_rsci_idat_3487_3456 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_0_sva, buf_linear_rsci_idat_3487_3456_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3519_3488 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_659 & (fsm_output[2]))
        | buf_linear_rsci_idat_3519_3488_mx0c1) ) begin
      buf_linear_rsci_idat_3519_3488 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_1_sva, buf_linear_rsci_idat_3519_3488_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3551_3520 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_659 & (fsm_output[2]))
        | buf_linear_rsci_idat_3551_3520_mx0c1) ) begin
      buf_linear_rsci_idat_3551_3520 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_2_sva, buf_linear_rsci_idat_3551_3520_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3583_3552 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_659 & (fsm_output[2]))
        | buf_linear_rsci_idat_3583_3552_mx0c1) ) begin
      buf_linear_rsci_idat_3583_3552 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_3_sva, buf_linear_rsci_idat_3583_3552_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3615_3584 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_677 & (fsm_output[2]))
        | buf_linear_rsci_idat_3615_3584_mx0c1) ) begin
      buf_linear_rsci_idat_3615_3584 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_4_sva, buf_linear_rsci_idat_3615_3584_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3647_3616 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_677 & (fsm_output[2]))
        | buf_linear_rsci_idat_3647_3616_mx0c1) ) begin
      buf_linear_rsci_idat_3647_3616 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_5_sva, buf_linear_rsci_idat_3647_3616_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3679_3648 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_677 & (fsm_output[2]))
        | buf_linear_rsci_idat_3679_3648_mx0c1) ) begin
      buf_linear_rsci_idat_3679_3648 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_6_sva, buf_linear_rsci_idat_3679_3648_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3711_3680 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_677 & (fsm_output[2]))
        | buf_linear_rsci_idat_3711_3680_mx0c1) ) begin
      buf_linear_rsci_idat_3711_3680 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_7_sva, buf_linear_rsci_idat_3711_3680_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3743_3712 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_694 & (fsm_output[2]))
        | buf_linear_rsci_idat_3743_3712_mx0c1) ) begin
      buf_linear_rsci_idat_3743_3712 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_8_sva, buf_linear_rsci_idat_3743_3712_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3775_3744 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_694 & (fsm_output[2]))
        | buf_linear_rsci_idat_3775_3744_mx0c1) ) begin
      buf_linear_rsci_idat_3775_3744 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_9_sva, buf_linear_rsci_idat_3775_3744_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3807_3776 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_694 & (fsm_output[2]))
        | buf_linear_rsci_idat_3807_3776_mx0c1) ) begin
      buf_linear_rsci_idat_3807_3776 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_10_sva, buf_linear_rsci_idat_3807_3776_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3839_3808 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_694 & (fsm_output[2]))
        | buf_linear_rsci_idat_3839_3808_mx0c1) ) begin
      buf_linear_rsci_idat_3839_3808 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_11_sva, buf_linear_rsci_idat_3839_3808_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3871_3840 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_711 & (fsm_output[2]))
        | buf_linear_rsci_idat_3871_3840_mx0c1) ) begin
      buf_linear_rsci_idat_3871_3840 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_12_sva, buf_linear_rsci_idat_3871_3840_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3903_3872 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_711 & (fsm_output[2]))
        | buf_linear_rsci_idat_3903_3872_mx0c1) ) begin
      buf_linear_rsci_idat_3903_3872 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_13_sva, buf_linear_rsci_idat_3903_3872_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3935_3904 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_194 & and_dcpl_711 & (fsm_output[2]))
        | buf_linear_rsci_idat_3935_3904_mx0c1) ) begin
      buf_linear_rsci_idat_3935_3904 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_14_sva, buf_linear_rsci_idat_3935_3904_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3967_3936 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_200 & and_dcpl_711 & (fsm_output[2]))
        | buf_linear_rsci_idat_3967_3936_mx0c1) ) begin
      buf_linear_rsci_idat_3967_3936 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_15_sva, buf_linear_rsci_idat_3967_3936_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_3999_3968 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_174 & and_dcpl_728 & (fsm_output[2]))
        | buf_linear_rsci_idat_3999_3968_mx0c1) ) begin
      buf_linear_rsci_idat_3999_3968 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_16_sva, buf_linear_rsci_idat_3999_3968_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      buf_linear_rsci_idat_4031_4000 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & ((and_dcpl_178 & and_dcpl_188 & and_dcpl_728 & (fsm_output[2]))
        | buf_linear_rsci_idat_4031_4000_mx0c1) ) begin
      buf_linear_rsci_idat_4031_4000 <= MUX_v_32_2_2(LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0,
          LOAD_BATCH_LOOP_buf_tmp_lin_data_6_17_sva, buf_linear_rsci_idat_4031_4000_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse
          <= 1'b0;
      reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse
          <= 1'b0;
      reg_done_rsci_ivld_core_psct_cse <= 1'b0;
      reg_dma_read_ctrl_rsci_ivld_core_psct_cse <= 1'b0;
      reg_conf_info_rsci_irdy_core_psct_cse <= 1'b0;
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d_reg <= 14'b00000000000000;
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d_reg <= 14'b00000000000000;
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d_reg <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen ) begin
      reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse
          <= and_2370_rmff;
      reg_LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse
          <= and_2372_rmff;
      reg_done_rsci_ivld_core_psct_cse <= and_dcpl_24 & (fsm_output[2]);
      reg_dma_read_ctrl_rsci_ivld_core_psct_cse <= (mux_310_nl | LOAD_LOOP_for_LOAD_LOOP_nand_cse)
          & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
      reg_conf_info_rsci_irdy_core_psct_cse <= ~((fsm_output[2:1]!=2'b00));
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d_reg <= LOAD_LOOP_for_if_2_for_for_if_index_in_mux_rmff;
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d_reg <= LOAD_LOOP_for_if_2_for_for_else_index_in_mux_rmff;
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d_reg <= LOAD_LOOP_for_if_2_for_for_if_mux_rmff;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_read_chnl_rsci_irdy_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((~((~ (fsm_output[2])) | mux_296_nl)) | or_tmp_2017) )
        begin
      reg_dma_read_chnl_rsci_irdy_core_psct_cse <= (~((~ mux_274_nl) & and_dcpl_738
          & (fsm_output[2]))) | or_tmp_2017;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_kernel_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_44 & (fsm_output[2])) | or_tmp_2027) ) begin
      reg_plm_kernel_rsci_ivld_core_psct_cse <= ~ or_tmp_2027;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_buf_linear_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_2033 | (or_tmp_4 & or_9_cse & and_dcpl_183 & (fsm_output[2])))
        ) begin
      reg_buf_linear_rsci_ivld_core_psct_cse <= ~ or_tmp_2033;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_asn_itm_2 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0 <= 2'b00;
      exitL_exit_LOAD_LOOP_for_if_2_for_sva_1 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2 <= 1'b0;
      LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3 <= 3'b000;
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4 <= 3'b000;
      sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1 <= 1'b0;
      LOAD_LOOP_for_print_buf_lpi_2_dfm_3 <= 8'b00000000;
      LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3 <= 5'b00000;
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4 <= 5'b00000;
    end
    else if ( LOAD_LOOP_for_if_for_and_cse ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_2 <= exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_1;
      LOAD_LOOP_for_if_2_for_for_asn_itm_2 <= LOAD_LOOP_for_if_2_for_for_asn_itm_1;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0;
      exitL_exit_LOAD_LOOP_for_if_2_for_sva_1 <= exitL_exit_LOAD_LOOP_for_if_2_for_sva_1_mx0w0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2_mx0w0;
      LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3 <= LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3_mx0w0;
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4 <= LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4_mx0w0;
      sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1 <= sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1_mx0w0;
      LOAD_LOOP_for_print_buf_lpi_2_dfm_3 <= LOAD_LOOP_for_print_buf_lpi_2_dfm_3_mx0w0;
      LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3 <= LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3_mx0w0;
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4 <= LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3 <= 1'b0;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0 <= 2'b00;
    end
    else if ( LOAD_LOOP_for_if_2_for_if_and_128_cse ) begin
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_3 <= LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_2;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_3 <= exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_2;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_2 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_3_1_0 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | and_3197_cse | mux_336_nl | or_dcpl_136))
        ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm <= exit_LOAD_LOOP_for_if_for_lpi_2_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | or_dcpl_147 | or_dcpl_146)) ) begin
      exit_LOAD_LOOP_lpi_2_dfm_1 <= exit_LOAD_LOOP_lpi_2_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm <= 1'b0;
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_2_for_and_205_cse ) begin
      exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm <= or_810_cse;
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st <= LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_equal_tmp_2_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_or_tmp_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_equal_tmp_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_nor_tmp_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_mux_11_itm_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_equal_tmp_1_1 <= 1'b0;
      exit_LOAD_LOOP_for_if_2_for_for_sva_1 <= 1'b0;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_1 <= 1'b0;
      exit_LOAD_LOOP_for_if_2_for_sva_1_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_1 <= 1'b0;
      LOAD_LOOP_for_asn_2_itm_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_asn_itm_1 <= 1'b0;
      LOAD_BATCH_LOOP_asn_itm_1 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0 <= 2'b00;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0
          <= 3'b000;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_5_3
          <= 3'b000;
      exit_LOAD_LOOP_for_lpi_2_dfm_3 <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_for_and_2_cse ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st_1 <= MUX_s_1_2_2(exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0,
          exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st, or_tmp_2056);
      LOAD_LOOP_for_if_2_for_equal_tmp_2_1 <= LOAD_LOOP_for_if_2_for_equal_tmp_2_mx0w0;
      LOAD_LOOP_for_if_2_for_or_tmp_1 <= LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_and_cse_1
          | LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_nor_1_cse_1;
      LOAD_LOOP_for_if_2_for_equal_tmp_1 <= LOAD_LOOP_for_if_2_for_equal_tmp_mx0w0;
      LOAD_LOOP_for_if_2_for_nor_tmp_1 <= ~(LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_and_cse_1
          | LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_nor_1_cse_1 | LOAD_LOOP_for_if_2_for_equal_tmp_mx0w0
          | LOAD_LOOP_for_if_2_for_equal_tmp_1_mx0w0 | LOAD_LOOP_for_if_2_for_equal_tmp_2_mx0w0);
      LOAD_LOOP_for_if_2_for_mux_11_itm_1 <= MUX_s_1_2_2(LOAD_LOOP_for_if_for_LOAD_LOOP_for_if_for_or_1_nl,
          sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_mx1, or_tmp_2056);
      LOAD_LOOP_for_if_2_for_equal_tmp_1_1 <= LOAD_LOOP_for_if_2_for_equal_tmp_1_mx0w0;
      exit_LOAD_LOOP_for_if_2_for_for_sva_1 <= LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_if_1_LOAD_LOOP_for_if_2_for_for_if_1_nor_tmp;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_1 <= exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0;
      exit_LOAD_LOOP_for_if_2_for_sva_1_1 <= LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_1_LOAD_LOOP_for_if_2_for_if_1_nor_tmp;
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_1 <= LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_mx0w0;
      LOAD_LOOP_for_asn_2_itm_1 <= MUX_s_1_2_2(LOAD_LOOP_for_asn_sft_lpi_2, LOAD_LOOP_for_asn_2_itm,
          and_2516_nl);
      LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st_1 <= MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_mx0w1,
          LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st, and_2526_nl);
      LOAD_LOOP_for_if_2_for_for_asn_itm_1 <= MUX_s_1_2_2(operator_8_false_operator_8_false_nor_cse_lpi_2,
          LOAD_LOOP_for_if_2_for_for_asn_itm, or_tmp_2094);
      LOAD_BATCH_LOOP_asn_itm_1 <= LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse
          & exit_LOAD_LOOP_lpi_2_dfm_4;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_1 <= MUX_s_1_2_2(exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0,
          exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st, and_2666_nl);
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0
          <= MUX_v_3_2_2((LOAD_LOOP_for_if_2_for_for_acc_2_psp_1[2:0]), LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_0,
          or_tmp_2094);
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_5_3
          <= MUX_v_3_2_2(LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3_mx0w0,
          LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3,
          or_tmp_2094);
      exit_LOAD_LOOP_for_lpi_2_dfm_3 <= exit_LOAD_LOOP_for_lpi_2_dfm_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1 <= 6'b000000;
    end
    else if ( core_wen & mux_390_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2])
        ) begin
      LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1 <= nl_LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_1_0 <= 2'b00;
    end
    else if ( core_wen & mux_393_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2])
        ) begin
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_1_0 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_0_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_1 <= 1'b0;
      LOAD_LOOP_for_if_for_for_n_2_0_sva_1_1 <= 3'b000;
      exit_LOAD_LOOP_for_if_for_for_sva_1 <= 1'b0;
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_2_1 <= 3'b000;
      exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_1 <= 1'b0;
      LOAD_LOOP_for_if_for_m_2_0_sva_1_1 <= 3'b000;
      exit_LOAD_LOOP_for_if_for_sva_1_1 <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_for_and_3_cse ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_1 <= exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0;
      LOAD_LOOP_for_if_for_for_n_2_0_sva_1_1 <= LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1;
      exit_LOAD_LOOP_for_if_for_for_sva_1 <= exit_LOAD_LOOP_for_if_for_for_sva_mx0w0;
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_2_1 <= MUX_v_3_2_2(3'b000, LOAD_LOOP_for_if_for_for_if_mux_nl,
          exit_LOAD_LOOP_for_if_for_lpi_2_dfm_mx0w0);
      exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_1 <= exit_LOAD_LOOP_for_if_for_for_lpi_2_dfm_mx0w0;
      LOAD_LOOP_for_if_for_m_2_0_sva_1_1 <= LOAD_LOOP_for_if_for_m_2_0_sva_1_mx0w1;
      exit_LOAD_LOOP_for_if_for_sva_1_1 <= exit_LOAD_LOOP_for_if_for_sva_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_1 <= 5'b00000;
    end
    else if ( core_wen & and_dcpl_778 & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2])
        ) begin
      LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_1 <= LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_2_1 <= 5'b00000;
      LOAD_LOOP_for_print_buf_sva_1_1 <= 8'b00000000;
      LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1 <= 14'b00000000000000;
      LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_1 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_2_for_for_col_and_2_cse ) begin
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_2_1 <= MUX_v_5_2_2(5'b00000, LOAD_LOOP_for_if_2_for_for_if_1_mux_nl,
          or_810_cse);
      LOAD_LOOP_for_print_buf_sva_1_1 <= nl_LOAD_LOOP_for_print_buf_sva_1_1[7:0];
      LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1 <= nl_LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1[13:0];
      LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_1 <= LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_mx0w1;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_4_1_2 <= ~ exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_row_4_0_sva_1_1 <= 5'b00000;
    end
    else if ( core_wen & (~ LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_1_LOAD_LOOP_for_if_2_for_if_1_nor_tmp)
        & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]) ) begin
      LOAD_LOOP_for_if_2_for_row_4_0_sva_1_1 <= LOAD_LOOP_for_if_2_for_row_4_0_sva_1_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_asn_6_itm_1 <= 1'b0;
    end
    else if ( core_wen & mux_409_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2])
        ) begin
      LOAD_LOOP_for_asn_6_itm_1 <= LOAD_LOOP_for_asn_sft_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2 <= 1'b0;
    end
    else if ( core_wen & mux_476_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2])
        ) begin
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_2_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_for_for_and_108_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_107_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_106_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_105_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_104_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_103_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_102_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_101_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_100_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_99_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_98_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_97_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_96_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_95_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_94_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_93_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_92_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_91_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_90_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_89_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_88_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_87_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_86_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_85_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_84_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_83_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_82_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_81_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_80_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_79_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_78_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_77_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_76_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_75_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_74_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_73_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_72_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_71_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_70_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_69_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_68_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_67_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_66_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_65_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_64_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_63_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_62_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_61_psp <= 1'b0;
      LOAD_LOOP_for_if_for_for_and_60_psp <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_for_for_and_111_cse ) begin
      LOAD_LOOP_for_if_for_for_and_108_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_16_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_107_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_0_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_106_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_15_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_105_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_1_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_104_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_14_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_103_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_2_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_102_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_13_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_101_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_3_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_100_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_12_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_99_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_4_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_98_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_11_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_97_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_5_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_96_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_10_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_95_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_6_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_94_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_9_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_93_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_7_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_92_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_8_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_91_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_8_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_90_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_7_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_89_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_9_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_88_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_6_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_87_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_10_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_86_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_5_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_85_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_11_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_84_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_4_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_83_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_12_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_82_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_3_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_81_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_13_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_80_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_2_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_79_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_14_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_78_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_1_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_77_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_15_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_76_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_0_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]);
      LOAD_LOOP_for_if_for_for_and_75_psp <= LOAD_LOOP_for_if_for_for_and_stg_4_16_sva_1
          & (~ (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5]));
      LOAD_LOOP_for_if_for_for_and_74_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_15_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_73_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_1_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_72_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_14_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_71_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_2_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_70_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_13_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_69_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_3_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_68_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_12_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_67_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_4_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_66_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_11_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_65_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_5_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_64_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_10_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_63_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_6_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_62_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_9_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_61_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_7_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
      LOAD_LOOP_for_if_for_for_and_60_psp <= LOAD_LOOP_for_if_for_for_and_stg_3_8_sva_1
          & (LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1[5:4]==2'b01);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_asn_2_itm <= 1'b0;
    end
    else if ( LOAD_LOOP_for_and_2_cse & (~(mux_481_cse | or_dcpl_136)) ) begin
      LOAD_LOOP_for_asn_2_itm <= LOAD_LOOP_for_asn_sft_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | mux_tmp_353 | LOAD_LOOP_for_LOAD_LOOP_nand_cse
        | (~(LOAD_BATCH_LOOP_and_4_tmp & operator_8_false_operator_8_false_nor_cse_lpi_2))))
        ) begin
      LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_st <= LOAD_LOOP_for_if_2_for_for_if_land_2_lpi_2_dfm_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_for_asn_itm <= 1'b0;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3
          <= 3'b000;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_0
          <= 3'b000;
    end
    else if ( LOAD_LOOP_for_if_2_for_for_and_257_cse ) begin
      LOAD_LOOP_for_if_2_for_for_asn_itm <= operator_8_false_operator_8_false_nor_cse_lpi_2;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st <= exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3
          <= LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_5_3_mx0w0;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_0
          <= LOAD_LOOP_for_if_2_for_for_acc_2_psp_1[2:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1 <= 1'b0;
    end
    else if ( core_wen & (((~ mux_515_nl) & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0
        & and_dcpl_752 & (fsm_output[2])) | LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1_mx0c1)
        ) begin
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1 <= MUX_s_1_2_2(LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_mx0w0,
          LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st, LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st <= 1'b0;
    end
    else if ( LOAD_LOOP_for_and_2_cse & (~(mux_tmp_575 | or_dcpl_136)) ) begin
      exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_st <= exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_for_and_249_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_248_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_247_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_246_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_245_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_244_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_243_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_242_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_241_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_240_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_239_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_238_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_237_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_236_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_235_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_234_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_233_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_232_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_231_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_230_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_229_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_228_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_227_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_226_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_225_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_224_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_223_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_222_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_221_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_220_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_219_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_218_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_217_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_216_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_215_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_214_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_213_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_212_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_211_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_210_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_209_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_208_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_207_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_206_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_205_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_204_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_203_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_202_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_201_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_200_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_199_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_198_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_197_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_196_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_195_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_194_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_193_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_192_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_191_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_190_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_189_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_188_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_187_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_186_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_185_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_184_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_183_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_182_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_181_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_180_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_179_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_178_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_177_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_176_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_175_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_174_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_173_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_172_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_171_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_170_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_169_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_168_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_167_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_166_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_165_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_164_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_163_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_162_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_161_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_160_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_159_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_158_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_157_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_156_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_155_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_154_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_153_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_152_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_151_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_150_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_149_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_148_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_147_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_146_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_145_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_144_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_143_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_142_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_141_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_140_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_139_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_138_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_137_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_136_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_135_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_134_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_133_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_132_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_131_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_130_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_129_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_128_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_127_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_126_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_125_psp <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_124_psp <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_2_for_for_and_259_cse ) begin
      LOAD_LOOP_for_if_2_for_for_and_249_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_61_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_248_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_0_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_247_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_60_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_246_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_1_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_245_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_59_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_244_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_2_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_243_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_58_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_242_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_3_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_241_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_57_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_240_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_4_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_239_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_56_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_238_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_5_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_237_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_55_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_236_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_6_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_235_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_54_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_234_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_7_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_233_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_53_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_232_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_8_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_231_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_52_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_230_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_9_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_229_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_51_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_228_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_10_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_227_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_50_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_226_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_11_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_225_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_49_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_224_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_12_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_223_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_48_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_222_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_13_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_221_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_47_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_220_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_14_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_219_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_46_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_218_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_15_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_217_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_45_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_216_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_16_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_215_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_44_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_214_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_17_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_213_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_43_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_212_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_18_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_211_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_42_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_210_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_19_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_209_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_41_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_208_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_20_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_207_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_40_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_206_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_21_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_205_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_39_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_204_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_22_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_203_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_38_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_202_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_23_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_201_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_37_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_200_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_24_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_199_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_36_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_198_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_25_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_197_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_35_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_196_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_26_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_195_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_34_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_194_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_27_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_193_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_33_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_192_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_28_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_191_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_32_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_190_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_29_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_189_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_31_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_188_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_30_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_187_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_30_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_186_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_31_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_185_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_29_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_184_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_32_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_183_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_28_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_182_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_33_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_181_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_27_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_180_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_34_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_179_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_26_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_178_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_35_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_177_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_25_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_176_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_36_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_175_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_24_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_174_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_37_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_173_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_23_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_172_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_38_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_171_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_22_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_170_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_39_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_169_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_21_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_168_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_40_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_167_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_20_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_166_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_41_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_165_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_19_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_164_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_42_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_163_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_18_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_162_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_43_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_161_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_17_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_160_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_44_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_159_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_16_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_158_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_45_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_157_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_15_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_156_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_46_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_155_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_14_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_154_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_47_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_153_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_13_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_152_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_48_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_151_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_12_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_150_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_49_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_149_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_11_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_148_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_50_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_147_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_10_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_146_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_51_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_145_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_9_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_144_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_52_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_143_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_8_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_142_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_53_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_141_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_7_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_140_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_54_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_139_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_6_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_138_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_55_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_137_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_5_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_136_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_56_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_135_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_4_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_134_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_57_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_133_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_3_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_132_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_58_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_131_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_2_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_130_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_59_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_129_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_1_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_128_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_60_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_127_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_0_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]);
      LOAD_LOOP_for_if_2_for_for_and_126_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_5_61_sva_1
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2]));
      LOAD_LOOP_for_if_2_for_for_and_125_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_4_31_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b01);
      LOAD_LOOP_for_if_2_for_for_and_124_psp <= LOAD_LOOP_for_if_2_for_for_and_stg_4_30_sva_1
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]==2'b01);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0 <= 2'b00;
    end
    else if ( core_wen & (~((fsm_output[3]) | (fsm_output[0]) | ((~ LOAD_BATCH_LOOP_and_3_tmp)
        & (fsm_output[2])))) ) begin
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0 <= lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1 <= 1'b0;
      LOAD_LOOP_for_asn_sft_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( operator_8_false_and_cse ) begin
      operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1 <= MUX_s_1_2_2(LOAD_LOOP_for_if_for_mux_11_nl,
          operator_8_false_operator_8_false_nor_cse_lpi_2, or_tmp_2315);
      LOAD_LOOP_for_asn_sft_lpi_2_dfm_1 <= MUX_s_1_2_2(LOAD_LOOP_for_if_for_mux_12_nl,
          LOAD_LOOP_for_asn_sft_lpi_2, or_tmp_2315);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2 <= 16'b0000000000000000;
    end
    else if ( core_wen & (or_tmp_1481 | LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2_mx0c1)
        ) begin
      LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2 <= MUX_v_16_2_2((z_out_10[15:0]),
          LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2, LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_v <= 1'b0;
    end
    else if ( core_wen & (LOAD_BATCH_LOOP_stage_v_mx0c0 | LOAD_BATCH_LOOP_stage_v_mx0c1)
        ) begin
      LOAD_BATCH_LOOP_stage_v <= (~ LOAD_BATCH_LOOP_stage_v_mx0c1) | LOAD_BATCH_LOOP_stage_v_mx0c0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (LOAD_BATCH_LOOP_stage_v_2_mx0c0 | (LOAD_BATCH_LOOP_and_3_tmp
        & (fsm_output[2]))) ) begin
      LOAD_BATCH_LOOP_stage_v_2 <= ~ LOAD_BATCH_LOOP_stage_v_2_mx0c0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_2 <= 1'b0;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_2 <= 1'b0;
      LOAD_BATCH_LOOP_asn_itm_2 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3
          <= 3'b000;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1
          <= 2'b00;
      LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 <= 1'b0;
      LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1 <= 32'b00000000000000000000000000000000;
      LOAD_LOOP_for_if_2_for_for_asn_126_itm_2 <= 1'b0;
      LOAD_LOOP_for_if_2_for_equal_tmp_2_2 <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_2_for_if_and_132_cse ) begin
      LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_2 <= LOAD_LOOP_for_if_2_for_LOAD_LOOP_for_if_2_for_if_and_svs_st_1;
      exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_2 <= exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_st_1;
      LOAD_BATCH_LOOP_asn_itm_2 <= LOAD_BATCH_LOOP_asn_itm_1;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3
          <= LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_5_3;
      LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1
          <= LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0[2:1];
      LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 <= (~ (LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2[0]))
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0[0]);
      LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 <= (LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2[0])
          & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0[0]);
      LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 <= ~((LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2[0])
          | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0[0]));
      LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 <= (LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2[0])
          & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_1_2_0[0]));
      LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1 <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_mx0w0;
      LOAD_LOOP_for_if_2_for_for_asn_126_itm_2 <= LOAD_LOOP_for_if_2_for_for_asn_itm_1;
      LOAD_LOOP_for_if_2_for_equal_tmp_2_2 <= LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (LOAD_BATCH_LOOP_stage_v_3_mx0c0 | (and_dcpl_831 & (fsm_output[2])))
        ) begin
      LOAD_BATCH_LOOP_stage_v_3 <= ~ LOAD_BATCH_LOOP_stage_v_3_mx0c0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2 <= 3'b000;
      LOAD_LOOP_for_if_for_m_2_0_lpi_2 <= 3'b000;
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2 <= 5'b00000;
      LOAD_LOOP_for_if_2_for_row_4_0_lpi_2 <= 5'b00000;
      sfi_operator_8_false_operator_8_false_nor_cse_lpi_2 <= 1'b0;
      LOAD_LOOP_for_print_buf_lpi_2 <= 8'b00000000;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0 <= 2'b00;
      exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 <= 1'b0;
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2 <= 1'b0;
    end
    else if ( LOAD_LOOP_for_if_for_for_n_and_1_cse ) begin
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2 <= MUX_v_3_2_2(LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4,
          LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_dfm_4_mx0w0, or_tmp_2337);
      LOAD_LOOP_for_if_for_m_2_0_lpi_2 <= MUX_v_3_2_2(LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3,
          LOAD_LOOP_for_if_for_m_2_0_lpi_2_dfm_3_mx0w0, or_tmp_2337);
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2 <= MUX_v_5_2_2(LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4,
          LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_dfm_4_mx0w0, or_tmp_2337);
      LOAD_LOOP_for_if_2_for_row_4_0_lpi_2 <= MUX_v_5_2_2(LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3,
          LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_dfm_3_mx0w0, or_tmp_2337);
      sfi_operator_8_false_operator_8_false_nor_cse_lpi_2 <= MUX_s_1_2_2(sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1,
          sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1_mx0w0, or_tmp_2337);
      LOAD_LOOP_for_print_buf_lpi_2 <= MUX_v_8_2_2(LOAD_LOOP_for_print_buf_lpi_2_dfm_3,
          LOAD_LOOP_for_print_buf_lpi_2_dfm_3_mx0w0, or_tmp_2337);
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0 <= MUX_v_2_2_2(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0,
          lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_1_0_mx0w0, or_tmp_2337);
      exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 <= MUX_s_1_2_2(exitL_exit_LOAD_LOOP_for_if_2_for_sva_1,
          exitL_exit_LOAD_LOOP_for_if_2_for_sva_1_mx0w0, or_tmp_2337);
      lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2 <= MUX_s_1_2_2(lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2,
          lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_5_2_mx0w0, or_tmp_2337);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_crt_sva_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      batch_size_mul_3_cse_sva <= 16'b0000000000000000;
      batch_size_mul_4_cse_sva <= 16'b0000000000000000;
      batch_size_sva <= 16'b0000000000000000;
      batch_size_mul_1_cse_sva <= 16'b0000000000000000;
      n_w_in_acc_psp_sva <= 7'b0000000;
      pad_sva <= 8'b00000000;
      n_h_in_acc_psp_sva <= 7'b0000000;
      batch_size_mul_2_cse_sva <= 16'b0000000000000000;
    end
    else if ( and_cse ) begin
      conf_info_crt_sva_231_0 <= conf_info_rsci_idat_mxwt;
      batch_size_mul_3_cse_sva <= z_out_2_15_0;
      batch_size_mul_4_cse_sva <= z_out_15_0;
      batch_size_sva <= z_out_12;
      batch_size_mul_1_cse_sva <= z_out_3_15_0;
      n_w_in_acc_psp_sva <= nl_n_w_in_acc_psp_sva[6:0];
      pad_sva <= z_out_1[7:0];
      n_h_in_acc_psp_sva <= nl_n_h_in_acc_psp_sva[6:0];
      batch_size_mul_2_cse_sva <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_0 <= 1'b0;
    end
    else if ( core_wen & ((fsm_output[1]) | or_tmp_2350) ) begin
      LOAD_BATCH_LOOP_stage_0 <= ~ or_tmp_2350;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_fl_5_0_sva_4_0 <= 5'b00000;
      lfst_exit_LOAD_LOOP_sva <= 1'b0;
      lfst_exit_LOAD_LOOP_for_1_lpi_2 <= 1'b0;
    end
    else if ( LOAD_LOOP_fl_and_cse ) begin
      LOAD_LOOP_fl_5_0_sva_4_0 <= LOAD_LOOP_for_mux_7_nl & ({{4{lfst_exit_LOAD_LOOP_sva_dfm_1_mx0w1}},
          lfst_exit_LOAD_LOOP_sva_dfm_1_mx0w1}) & (signext_5_1(~ (fsm_output[1])));
      lfst_exit_LOAD_LOOP_sva <= lfst_exit_LOAD_LOOP_sva_dfm_1_mx0w1 & (~ (fsm_output[1]));
      lfst_exit_LOAD_LOOP_for_1_lpi_2 <= MUX_s_1_2_2((~ exit_LOAD_LOOP_for_lpi_2_dfm_3),
          (~ exit_LOAD_LOOP_for_lpi_2_dfm_3_mx0w0), or_tmp_2354);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_b_4_0_sva_3_0 <= 4'b0000;
    end
    else if ( core_wen & ((fsm_output[1]) | ((~ mux_tmp_597) & or_810_cse & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0
        & and_3266_cse & (~ LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_nor_tmp)
        & (~ (LOAD_BATCH_LOOP_acc_tmp[4])) & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2])))
        ) begin
      LOAD_BATCH_LOOP_b_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, (LOAD_BATCH_LOOP_acc_tmp[3:0]),
          LOAD_BATCH_LOOP_b_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_ac_int_cctor_lpi_2 <= 16'b0000000000000000;
      LOAD_LOOP_for_mul_cse_lpi_2 <= 16'b0000000000000000;
    end
    else if ( LOAD_LOOP_for_and_5_cse ) begin
      LOAD_LOOP_for_ac_int_cctor_lpi_2 <= z_out_10[15:0];
      LOAD_LOOP_for_mul_cse_lpi_2 <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2 <= 16'b0000000000000000;
    end
    else if ( core_wen & ((fsm_output[1]) | or_tmp_1481) ) begin
      LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2 <= MUX_v_16_2_2(LOAD_LOOP_for_if_1_ac_int_cctor_lpi_2_dfm_2,
          (z_out_10[15:0]), or_tmp_1481);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_asn_sft_lpi_2 <= 1'b0;
      operator_8_false_operator_8_false_nor_cse_lpi_2 <= 1'b0;
    end
    else if ( LOAD_LOOP_for_and_9_cse ) begin
      LOAD_LOOP_for_asn_sft_lpi_2 <= MUX_s_1_2_2(LOAD_LOOP_for_asn_sft_lpi_2_dfm_1,
          operator_8_false_operator_8_false_nor_cse_sva_1, or_tmp_2314);
      operator_8_false_operator_8_false_nor_cse_lpi_2 <= MUX_s_1_2_2(operator_8_false_operator_8_false_nor_cse_lpi_2_dfm_1,
          operator_8_false_operator_8_false_nor_cse_sva_1, or_tmp_2314);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_for_k_5_0_lpi_2_4_0 <= 5'b00000;
    end
    else if ( core_wen & (((~ mux_621_nl) & or_810_cse & exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0
        & (~ (LOAD_LOOP_acc_tmp[5])) & lfst_exit_LOAD_LOOP_for_1_lpi_2 & lfst_exit_LOAD_LOOP_sva
        & LOAD_BATCH_LOOP_and_4_tmp) | LOAD_LOOP_for_k_5_0_lpi_2_4_0_mx0c1) ) begin
      LOAD_LOOP_for_k_5_0_lpi_2_4_0 <= MUX1HOT_v_5_3_2(({{4{exit_LOAD_LOOP_lpi_2_dfm_1_mx0w0}},
          exit_LOAD_LOOP_lpi_2_dfm_1_mx0w0}), (LOAD_LOOP_for_acc_2_tmp[4:0]), LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1,
          {(~ LOAD_LOOP_for_k_5_0_lpi_2_4_0_mx0c1) , LOAD_LOOP_for_k_and_nl , LOAD_LOOP_for_k_and_1_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (LOAD_BATCH_LOOP_stage_v_1_mx0c0 | and_3158_cse) ) begin
      LOAD_BATCH_LOOP_stage_v_1 <= ~ LOAD_BATCH_LOOP_stage_v_1_mx0c0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_48_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_623_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_48_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_625_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_0_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_47_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_627_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_47_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_629_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_1_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_46_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_631_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_46_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_633_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_2_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_45_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_635_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_45_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_637_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_3_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_44_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_639_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_44_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_641_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_4_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_43_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_643_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_43_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_645_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_5_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_42_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_647_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_42_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_649_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_6_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_41_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_651_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_41_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_653_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_7_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_40_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_655_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_40_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_657_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_8_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_39_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_659_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_39_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_661_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_9_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_38_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_663_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_38_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_665_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_10_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_37_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_667_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_37_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_669_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_11_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_36_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_671_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_36_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_673_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_12_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_35_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_675_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_35_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_677_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_13_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_34_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_679_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_34_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_681_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_14_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_33_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_683_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_33_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_685_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_15_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_32_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_687_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_32_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_689_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_16_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_31_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_691_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_31_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_693_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_17_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_30_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_695_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_30_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_18_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_697_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_18_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_29_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_699_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_29_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_19_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_701_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_19_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_28_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_703_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_28_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_20_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_705_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_20_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_27_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_707_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_27_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_21_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_709_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_21_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_26_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_711_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_26_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_22_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_713_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_22_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_25_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_715_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_25_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_23_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_717_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_23_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_24_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~(mux_719_nl | or_dcpl_209)) ) begin
      LOAD_BATCH_LOOP_plm_tmp_f_data_24_sva <= dma_read_chnl_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_0_1 <= 1'b0;
    end
    else if ( core_wen & ((fsm_output[1]) | or_tmp_2350 | or_tmp_2354) ) begin
      LOAD_BATCH_LOOP_stage_0_1 <= (LOAD_BATCH_LOOP_stage_0 & (~ or_tmp_2350)) |
          (fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_0_2 <= 1'b0;
    end
    else if ( core_wen & ((fsm_output[1]) | ((LOAD_BATCH_LOOP_and_3_tmp | LOAD_BATCH_LOOP_and_4_tmp)
        & (fsm_output[2]))) ) begin
      LOAD_BATCH_LOOP_stage_0_2 <= LOAD_BATCH_LOOP_stage_0_1 & (~ (fsm_output[1]));
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_stage_0_3 <= 1'b0;
    end
    else if ( core_wen & ((fsm_output[1]) | ((and_dcpl_831 | LOAD_BATCH_LOOP_and_3_tmp)
        & (fsm_output[2]))) ) begin
      LOAD_BATCH_LOOP_stage_0_3 <= LOAD_BATCH_LOOP_stage_0_2 & (~ (fsm_output[1]));
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_722_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_17_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_725_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_0_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_728_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_16_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_731_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_1_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_734_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_15_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_737_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_2_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_740_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_14_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_743_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_3_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_746_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_13_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_749_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_4_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_752_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_12_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_755_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_5_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_758_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_11_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_761_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_6_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_764_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_10_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_767_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_7_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_770_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_9_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_773_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_8_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_776_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_8_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_779_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_9_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_782_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_7_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_785_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_10_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_788_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_6_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_791_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_11_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_794_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_5_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_797_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_12_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_800_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_4_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_803_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_13_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_806_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_3_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_809_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_14_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_812_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_2_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_815_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_15_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_818_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_1_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_821_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_16_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_824_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_6_0_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_827_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_0_17_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_830_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_17_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_833_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_0_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_836_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_16_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_839_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_1_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_842_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_15_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_845_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_2_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_848_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_14_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_851_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_3_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_854_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_13_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_857_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_4_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_860_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_12_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_863_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_5_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_866_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_11_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_869_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_6_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_872_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_10_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_875_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_7_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_878_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_9_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_881_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_8_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_884_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_8_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_887_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_9_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_890_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_7_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_893_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_10_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_896_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_6_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_899_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_11_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_902_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_5_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_905_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_12_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_908_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_4_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_911_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_13_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_914_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_3_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_917_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_14_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_920_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_2_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_923_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_15_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_926_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_1_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_929_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_16_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_932_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_5_0_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_935_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_1_17_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_938_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_17_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_941_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_0_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_944_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_16_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_947_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_1_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_950_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_15_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_953_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_2_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_956_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_14_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_959_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_3_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_962_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_13_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_965_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_4_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_968_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_12_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_971_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_5_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_974_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_11_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_977_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_6_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_980_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_10_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_983_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_7_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_986_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_9_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_989_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_8_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_992_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_8_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_995_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_9_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_998_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_7_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1001_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_10_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1004_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_6_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1007_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_11_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1010_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_5_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1013_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_12_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1016_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_4_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1019_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_13_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1022_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_3_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1025_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_14_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1028_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_2_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1031_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_15_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1034_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_1_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1037_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_16_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1040_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_4_0_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1043_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_2_17_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_17_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1046_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_17_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_0_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1049_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_0_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_16_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1052_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_16_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_1_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1055_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_1_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_15_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1058_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_15_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_2_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1061_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_2_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_14_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1064_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_14_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_3_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1067_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_3_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_13_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1070_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_13_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_4_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1073_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_4_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_12_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1076_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_12_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_5_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1079_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_5_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_11_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1082_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_11_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_6_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1085_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_6_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_10_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1088_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_10_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_7_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1091_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_7_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_9_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1094_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_9_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_8_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ mux_1097_nl) | or_dcpl_263)) ) begin
      LOAD_BATCH_LOOP_buf_tmp_lin_data_3_8_sva <= LOAD_LOOP_for_if_2_for_for_data_lpi_2_dfm_1_mx0;
    end
  end
  assign LOAD_CTRL_LOOP1_or_nl = ((~ and_1304_tmp) & or_tmp_1480) | or_tmp_1481;
  assign LOAD_CTRL_LOOP1_and_2_nl = and_1304_tmp & or_tmp_1480;
  assign or_485_nl = nor_tmp_67 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1]) | or_197_cse;
  assign or_483_nl = nor_tmp_63 | or_197_cse;
  assign mux_307_nl = MUX_s_1_2_2(or_485_nl, or_483_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_304_nl = MUX_s_1_2_2(nand_24_cse, mux_tmp_109, or_481_cse);
  assign mux_305_nl = MUX_s_1_2_2(mux_304_nl, nand_24_cse, nor_tmp_67);
  assign mux_303_nl = MUX_s_1_2_2(mux_tmp_109, nand_24_cse, nor_tmp_63);
  assign mux_306_nl = MUX_s_1_2_2(mux_305_nl, mux_303_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_308_nl = MUX_s_1_2_2(mux_307_nl, mux_306_nl, LOAD_LOOP_for_asn_sft_lpi_2);
  assign mux_309_nl = MUX_s_1_2_2(mux_107_cse, (~ mux_308_nl), LOAD_BATCH_LOOP_and_3_tmp);
  assign mux_310_nl = MUX_s_1_2_2(mux_309_nl, mux_107_cse, LOAD_BATCH_LOOP_asn_itm_1);
  assign mux_268_nl = MUX_s_1_2_2(nand_tmp_29, mux_tmp_260, or_481_cse);
  assign mux_267_nl = MUX_s_1_2_2(nand_tmp_29, mux_tmp_260, or_631_cse);
  assign mux_269_nl = MUX_s_1_2_2(mux_268_nl, mux_267_nl, nor_tmp_67);
  assign mux_266_nl = MUX_s_1_2_2(mux_tmp_260, nand_tmp_29, nor_tmp_63);
  assign mux_270_nl = MUX_s_1_2_2(mux_269_nl, mux_266_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_271_nl = MUX_s_1_2_2(mux_270_nl, nand_tmp_29, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign or_2861_nl = (~((lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b10) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2))
      | mux_tmp_260;
  assign or_2862_nl = (~((lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0!=2'b00) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2))
      | mux_tmp_260;
  assign mux_265_nl = MUX_s_1_2_2(or_2861_nl, or_2862_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2);
  assign mux_272_nl = MUX_s_1_2_2(mux_271_nl, mux_265_nl, LOAD_BATCH_LOOP_asn_itm_1);
  assign or_452_nl = nor_tmp_67 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b10);
  assign mux_262_nl = MUX_s_1_2_2(nand_tmp_29, mux_tmp_260, or_452_nl);
  assign or_451_nl = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 | LOAD_LOOP_for_if_2_for_equal_tmp_2_1;
  assign mux_263_nl = MUX_s_1_2_2(mux_262_nl, mux_tmp_260, or_451_nl);
  assign or_2868_nl = nor_778_cse | mux_tmp_260;
  assign mux_264_nl = MUX_s_1_2_2(mux_263_nl, or_2868_nl, LOAD_BATCH_LOOP_asn_itm_1);
  assign mux_273_nl = MUX_s_1_2_2(mux_272_nl, mux_264_nl, or_439_cse);
  assign mux_274_nl = MUX_s_1_2_2(mux_tmp_260, mux_273_nl, nor_tmp_101);
  assign or_474_nl = (~ LOAD_BATCH_LOOP_and_3_tmp) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0])
      | mux_tmp_260;
  assign mux_292_nl = MUX_s_1_2_2(nand_tmp_34, (~ or_tmp_352), lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1]);
  assign mux_291_nl = MUX_s_1_2_2((~ or_tmp_352), nand_tmp_34, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1]);
  assign mux_293_nl = MUX_s_1_2_2(mux_292_nl, mux_291_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2);
  assign or_467_nl = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[0]) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2;
  assign mux_294_nl = MUX_s_1_2_2(mux_293_nl, nand_tmp_34, or_467_nl);
  assign mux_281_nl = MUX_s_1_2_2(mux_1159_itm, or_tmp_340, or_461_itm);
  assign nor_725_nl = ~(or_75_cse | (~ mux_281_nl));
  assign mux_283_nl = MUX_s_1_2_2(nand_tmp_32, nor_725_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[1]);
  assign or_458_nl = (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_1_0[0]) | exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2
      | lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2;
  assign mux_284_nl = MUX_s_1_2_2(mux_283_nl, nand_tmp_32, or_458_nl);
  assign mux_295_nl = MUX_s_1_2_2(mux_294_nl, mux_284_nl, or_439_cse);
  assign mux_296_nl = MUX_s_1_2_2(or_474_nl, mux_295_nl, nor_tmp_101);
  assign or_538_nl = (~ or_tmp_154) | LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b10)
      | LOAD_LOOP_for_if_2_for_and_195_ssc_1 | and_834_cse;
  assign mux_336_nl = MUX_s_1_2_2(or_539_cse, or_538_nl, nor_37_cse);
  assign LOAD_LOOP_for_if_for_LOAD_LOOP_for_if_for_or_1_nl = sfi_operator_8_false_operator_8_false_nor_cse_lpi_2_mx1
      | exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0;
  assign nor_569_nl = ~((~((LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00))) | and_tmp_12);
  assign nor_571_nl = ~(((LOAD_LOOP_for_if_2_for_mux1h_378_tmp==2'b11)) | and_tmp_12);
  assign mux_421_nl = MUX_s_1_2_2(nor_569_nl, nor_571_nl, or_tmp_154);
  assign and_3194_nl = or_tmp_388 & (~ and_tmp_12);
  assign mux_422_nl = MUX_s_1_2_2(mux_421_nl, and_3194_nl, LOAD_LOOP_for_if_2_for_equal_tmp_2_1);
  assign mux_423_nl = MUX_s_1_2_2(mux_422_nl, and_tmp_12, LOAD_LOOP_for_if_2_for_and_195_ssc_1);
  assign mux_420_nl = MUX_s_1_2_2(not_tmp_236, or_632_cse, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_2);
  assign or_690_nl = exitL_exit_LOAD_LOOP_for_if_2_for_lpi_2 | mux_420_nl;
  assign mux_424_nl = MUX_s_1_2_2(mux_423_nl, or_690_nl, or_75_cse);
  assign mux_425_nl = MUX_s_1_2_2(mux_tmp_418, mux_424_nl, or_2860_cse);
  assign mux_426_nl = MUX_s_1_2_2(mux_tmp_418, mux_425_nl, or_513_cse);
  assign nand_55_nl = ~(and_3266_cse & (~ mux_426_nl));
  assign mux_427_nl = MUX_s_1_2_2(nand_tmp_52, nand_55_nl, LOAD_BATCH_LOOP_if_LOAD_BATCH_LOOP_if_or_1_cse);
  assign mux_428_nl = MUX_s_1_2_2(mux_427_nl, nand_tmp_52, nor_32_cse);
  assign mux_429_nl = MUX_s_1_2_2(nand_tmp_52, mux_428_nl, exit_LOAD_LOOP_for_if_2_for_for_lpi_2_dfm_mx0w0);
  assign and_872_nl = LOAD_BATCH_LOOP_stage_0 & mux_429_nl;
  assign mux_430_nl = MUX_s_1_2_2(and_872_nl, nand_tmp_52, or_588_cse);
  assign and_2516_nl = mux_430_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign nand_63_nl = ~(nor_tmp_172 & (~(nor_566_cse | LOAD_BATCH_LOOP_stage_0_3
      | LOAD_BATCH_LOOP_stage_0_2 | (LOAD_BATCH_LOOP_stage_0 & nand_tmp_62))));
  assign mux_468_nl = MUX_s_1_2_2(nand_63_nl, mux_tmp_457, operator_8_false_operator_8_false_nor_cse_lpi_2);
  assign and_2526_nl = mux_468_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign and_899_nl = LOAD_BATCH_LOOP_stage_0 & mux_tmp_456;
  assign mux_569_nl = MUX_s_1_2_2(mux_tmp_522, mux_tmp_456, LOAD_BATCH_LOOP_stage_0);
  assign mux_570_nl = MUX_s_1_2_2(and_899_nl, mux_569_nl, LOAD_BATCH_LOOP_stage_0_2);
  assign mux_571_nl = MUX_s_1_2_2(mux_570_nl, mux_tmp_456, or_771_cse);
  assign mux_572_nl = MUX_s_1_2_2(mux_571_nl, mux_tmp_456, LOAD_BATCH_LOOP_stage_0_1);
  assign and_2666_nl = mux_572_nl & LOAD_BATCH_LOOP_and_4_tmp & (fsm_output[2]);
  assign nl_LOAD_LOOP_for_if_for_for_index_f_acc_decb_sva_1  = (z_out_3_15_0[5:0])
      + conv_u2u_3_6(LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_mx1);
  assign nor_574_nl = ~((~((~ LOAD_LOOP_for_if_2_for_equal_tmp_1_1) | (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0[0])))
      | LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (~((LOAD_LOOP_for_if_2_for_mux1h_378_tmp[1])
      & or_tmp_471)));
  assign mux_389_nl = MUX_s_1_2_2(and_tmp_30, nor_574_nl, LOAD_BATCH_LOOP_and_3_tmp);
  assign mux_390_nl = MUX_s_1_2_2(mux_389_nl, and_tmp_30, LOAD_BATCH_LOOP_asn_itm_1);
  assign and_847_nl = or_632_cse & or_tmp_471;
  assign mux_391_nl = MUX_s_1_2_2(and_tmp_32, or_tmp_471, or_631_cse);
  assign and_3196_nl = LOAD_LOOP_for_if_2_for_equal_tmp_1_1 & (lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_1_0==2'b11)
      & (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_1_2) & dma_read_ctrl_rsci_irdy_mxwt
      & LOAD_LOOP_for_asn_2_itm_1;
  assign mux_392_nl = MUX_s_1_2_2(mux_391_nl, and_tmp_32, and_3196_nl);
  assign mux_393_nl = MUX_s_1_2_2(and_847_nl, mux_392_nl, nor_37_cse);
  assign LOAD_LOOP_for_if_for_for_if_mux_nl = MUX_v_3_2_2(LOAD_LOOP_for_if_for_for_n_2_0_sva_1_mx0w1,
      LOAD_LOOP_for_if_for_for_n_2_0_lpi_2_mx1, exit_LOAD_LOOP_for_if_for_for_sva_mx0w0);
  assign LOAD_LOOP_for_if_2_for_for_if_1_mux_nl = MUX_v_5_2_2(LOAD_LOOP_for_if_2_for_for_col_4_0_sva_1_mx0w1,
      LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1, LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_if_1_LOAD_LOOP_for_if_2_for_for_if_1_nor_tmp);
  assign nl_LOAD_LOOP_for_print_buf_sva_1_1  = conv_u2u_5_8(LOAD_LOOP_for_print_buf_lpi_2_mx1_4_0)
      + (conf_info_crt_sva_231_0[7:0]);
  assign LOAD_LOOP_for_if_2_for_for_if_index_in_mul_7_nl = conv_u2u_13_13(LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1
      * ({n_w_in_acc_psp_sva , (conf_info_crt_sva_231_0[192])}));
  assign nl_LOAD_LOOP_for_if_2_for_for_if_index_in_acc_3_nl = LOAD_LOOP_for_if_2_for_for_if_index_in_mul_7_nl
      + conv_u2u_5_13(LOAD_LOOP_for_if_2_for_for_col_4_0_lpi_2_mx1);
  assign LOAD_LOOP_for_if_2_for_for_if_index_in_acc_3_nl = nl_LOAD_LOOP_for_if_2_for_for_if_index_in_acc_3_nl[12:0];
  assign nl_LOAD_LOOP_for_if_2_for_for_if_index_in_acc_itm_1  = conv_u2u_13_14(LOAD_LOOP_for_if_2_for_for_if_index_in_acc_3_nl)
      + z_out_1;
  assign nand_48_nl = ~(LOAD_LOOP_for_if_2_for_and_195_ssc_1 & (~ mux_tmp_405));
  assign mux_407_nl = MUX_s_1_2_2(nand_48_nl, mux_tmp_405, nor_178_cse);
  assign mux_408_nl = MUX_s_1_2_2(and_tmp_30, (~ mux_407_nl), LOAD_BATCH_LOOP_and_3_tmp);
  assign mux_409_nl = MUX_s_1_2_2(mux_408_nl, and_tmp_30, LOAD_BATCH_LOOP_asn_itm_1);
  assign and_885_nl = or_755_cse & or_tmp_471;
  assign mux_471_nl = MUX_s_1_2_2(or_tmp_471, and_tmp_32, and_3192_cse);
  assign mux_470_nl = MUX_s_1_2_2(or_tmp_471, and_tmp_32, nor_225_cse);
  assign mux_472_nl = MUX_s_1_2_2(mux_471_nl, mux_470_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_469_nl = MUX_s_1_2_2(or_tmp_471, and_tmp_32, LOAD_LOOP_for_if_2_for_equal_tmp_1_1);
  assign mux_473_nl = MUX_s_1_2_2(mux_472_nl, mux_469_nl, or_750_cse);
  assign or_749_nl = LOAD_LOOP_for_if_2_for_equal_tmp_2_1 | (~ lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_1_2)
      | LOAD_LOOP_for_if_2_for_or_tmp_1 | (LOAD_LOOP_for_if_2_for_mux1h_378_tmp!=2'b00);
  assign mux_474_nl = MUX_s_1_2_2(and_tmp_32, mux_473_nl, or_749_nl);
  assign mux_475_nl = MUX_s_1_2_2(and_885_nl, mux_474_nl, nor_37_cse);
  assign mux_476_nl = MUX_s_1_2_2(or_tmp_471, mux_475_nl, and_3266_cse);
  assign mux_507_nl = MUX_s_1_2_2(mux_tmp_505, mux_tmp_502, nor_tmp_54);
  assign mux_509_nl = MUX_s_1_2_2(mux_510_cse, mux_507_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_511_nl = MUX_s_1_2_2(mux_510_cse, mux_509_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_512_nl = MUX_s_1_2_2(mux_510_cse, mux_511_nl, nor_752_cse);
  assign nand_69_nl = ~(LOAD_BATCH_LOOP_stage_0 & (~ mux_512_nl));
  assign mux_494_nl = MUX_s_1_2_2(nand_tmp_66, nand_tmp_65, nor_tmp_54);
  assign mux_496_nl = MUX_s_1_2_2(mux_497_cse, mux_494_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_498_nl = MUX_s_1_2_2(mux_497_cse, mux_496_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_499_nl = MUX_s_1_2_2(mux_497_cse, mux_498_nl, nor_752_cse);
  assign mux_488_nl = MUX_s_1_2_2(mux_tmp_486, mux_tmp_484, nor_tmp_54);
  assign mux_490_nl = MUX_s_1_2_2(mux_491_cse, mux_488_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_492_nl = MUX_s_1_2_2(mux_491_cse, mux_490_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_493_nl = MUX_s_1_2_2(mux_491_cse, mux_492_nl, nor_752_cse);
  assign mux_500_nl = MUX_s_1_2_2(mux_499_nl, mux_493_nl, LOAD_BATCH_LOOP_stage_0);
  assign mux_513_nl = MUX_s_1_2_2(nand_69_nl, mux_500_nl, LOAD_BATCH_LOOP_stage_0_2);
  assign mux_514_nl = MUX_s_1_2_2(mux_513_nl, mux_tmp_353, or_771_cse);
  assign mux_515_nl = MUX_s_1_2_2(mux_514_nl, mux_tmp_353, LOAD_BATCH_LOOP_stage_0_1);
  assign LOAD_LOOP_for_if_for_mux_11_nl = MUX_s_1_2_2(operator_8_false_operator_8_false_nor_cse_lpi_2,
      operator_8_false_operator_8_false_nor_cse_sva_1, exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0);
  assign LOAD_LOOP_for_if_for_mux_12_nl = MUX_s_1_2_2(LOAD_LOOP_for_asn_sft_lpi_2,
      operator_8_false_operator_8_false_nor_cse_sva_1, exit_LOAD_LOOP_for_if_for_lpi_2_dfm_2_mx0w0);
  assign nl_n_w_in_acc_psp_sva  = (conf_info_rsci_idat_mxwt[199:193]) + (z_out_1[6:0]);
  assign nl_n_h_in_acc_psp_sva  = (conf_info_rsci_idat_mxwt[167:161]) + (z_out_1[6:0]);
  assign LOAD_LOOP_for_and_1_nl = (~ exit_LOAD_LOOP_sva_3) & exit_LOAD_LOOP_for_lpi_2_dfm_3_mx0w0;
  assign LOAD_LOOP_for_mux_7_nl = MUX_v_5_2_2(LOAD_LOOP_fl_5_0_sva_4_0, (LOAD_LOOP_acc_tmp[4:0]),
      LOAD_LOOP_for_and_1_nl);
  assign LOAD_BATCH_LOOP_b_not_1_nl = ~ (fsm_output[1]);
  assign LOAD_LOOP_for_k_and_nl = (~ or_1873_tmp) & LOAD_LOOP_for_k_5_0_lpi_2_4_0_mx0c1;
  assign LOAD_LOOP_for_k_and_1_nl = or_1873_tmp & LOAD_LOOP_for_k_5_0_lpi_2_4_0_mx0c1;
  assign mux_616_nl = MUX_s_1_2_2(mux_tmp_614, mux_tmp_612, nor_tmp_54);
  assign mux_618_nl = MUX_s_1_2_2(mux_619_cse, mux_616_nl, LOAD_LOOP_for_asn_2_itm_1);
  assign mux_620_nl = MUX_s_1_2_2(mux_619_cse, mux_618_nl, LOAD_LOOP_for_asn_6_itm_1);
  assign mux_621_nl = MUX_s_1_2_2(mux_619_cse, mux_620_nl, nor_752_cse);
  assign mux_622_nl = MUX_s_1_2_2(or_dcpl_103, (~ LOAD_LOOP_for_if_for_for_and_108_psp),
      or_941_cse);
  assign nand_269_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_108_psp);
  assign mux_623_nl = MUX_s_1_2_2(mux_622_nl, nand_269_nl, or_939_cse);
  assign mux_624_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_107_psp),
      or_941_cse);
  assign nand_337_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_107_psp);
  assign mux_625_nl = MUX_s_1_2_2(mux_624_nl, nand_337_nl, or_939_cse);
  assign nand_336_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_106_psp);
  assign mux_626_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_106_psp),
      or_941_cse);
  assign mux_627_nl = MUX_s_1_2_2(nand_336_nl, mux_626_nl, and_3220_cse);
  assign mux_628_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_105_psp),
      or_941_cse);
  assign nand_268_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_105_psp);
  assign mux_629_nl = MUX_s_1_2_2(mux_628_nl, nand_268_nl, or_950_cse);
  assign nand_267_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_104_psp);
  assign mux_630_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_104_psp),
      or_941_cse);
  assign mux_631_nl = MUX_s_1_2_2(nand_267_nl, mux_630_nl, nor_302_cse);
  assign nand_266_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_103_psp);
  assign mux_632_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_103_psp),
      or_941_cse);
  assign mux_633_nl = MUX_s_1_2_2(nand_266_nl, mux_632_nl, nor_304_cse);
  assign mux_634_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_102_psp),
      or_941_cse);
  assign nand_265_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_102_psp);
  assign mux_635_nl = MUX_s_1_2_2(mux_634_nl, nand_265_nl, or_960_cse);
  assign nand_264_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_101_psp);
  assign mux_636_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_101_psp),
      or_941_cse);
  assign mux_637_nl = MUX_s_1_2_2(nand_264_nl, mux_636_nl, nor_307_cse);
  assign mux_638_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_100_psp),
      or_941_cse);
  assign nand_263_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_100_psp);
  assign mux_639_nl = MUX_s_1_2_2(mux_638_nl, nand_263_nl, or_967_cse);
  assign mux_640_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_99_psp),
      or_941_cse);
  assign nand_262_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_99_psp);
  assign mux_641_nl = MUX_s_1_2_2(mux_640_nl, nand_262_nl, or_967_cse);
  assign nand_261_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_98_psp);
  assign mux_642_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_98_psp),
      or_941_cse);
  assign mux_643_nl = MUX_s_1_2_2(nand_261_nl, mux_642_nl, nor_307_cse);
  assign mux_644_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_97_psp),
      or_941_cse);
  assign nand_260_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_97_psp);
  assign mux_645_nl = MUX_s_1_2_2(mux_644_nl, nand_260_nl, or_960_cse);
  assign nand_259_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_96_psp);
  assign mux_646_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_96_psp),
      or_941_cse);
  assign mux_647_nl = MUX_s_1_2_2(nand_259_nl, mux_646_nl, nor_304_cse);
  assign nand_258_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_95_psp);
  assign mux_648_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_95_psp),
      or_941_cse);
  assign mux_649_nl = MUX_s_1_2_2(nand_258_nl, mux_648_nl, nor_302_cse);
  assign mux_650_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_94_psp),
      or_941_cse);
  assign nand_257_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_94_psp);
  assign mux_651_nl = MUX_s_1_2_2(mux_650_nl, nand_257_nl, or_950_cse);
  assign nand_256_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_93_psp);
  assign mux_652_nl = MUX_s_1_2_2(or_dcpl_32, (~ LOAD_LOOP_for_if_for_for_and_93_psp),
      or_941_cse);
  assign mux_653_nl = MUX_s_1_2_2(nand_256_nl, mux_652_nl, and_3220_cse);
  assign mux_654_nl = MUX_s_1_2_2(or_dcpl_94, (~ LOAD_LOOP_for_if_for_for_and_92_psp),
      or_941_cse);
  assign nand_255_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_92_psp);
  assign mux_655_nl = MUX_s_1_2_2(mux_654_nl, nand_255_nl, or_939_cse);
  assign mux_656_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_91_psp),
      or_941_cse);
  assign nand_335_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_91_psp);
  assign mux_657_nl = MUX_s_1_2_2(mux_656_nl, nand_335_nl, or_939_cse);
  assign nand_334_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_90_psp);
  assign mux_658_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_90_psp),
      or_941_cse);
  assign mux_659_nl = MUX_s_1_2_2(nand_334_nl, mux_658_nl, and_3220_cse);
  assign mux_660_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_89_psp),
      or_941_cse);
  assign nand_254_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_89_psp);
  assign mux_661_nl = MUX_s_1_2_2(mux_660_nl, nand_254_nl, or_950_cse);
  assign nand_253_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_88_psp);
  assign mux_662_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_88_psp),
      or_941_cse);
  assign mux_663_nl = MUX_s_1_2_2(nand_253_nl, mux_662_nl, nor_302_cse);
  assign nand_252_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_87_psp);
  assign mux_664_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_87_psp),
      or_941_cse);
  assign mux_665_nl = MUX_s_1_2_2(nand_252_nl, mux_664_nl, nor_304_cse);
  assign mux_666_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_86_psp),
      or_941_cse);
  assign nand_251_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_86_psp);
  assign mux_667_nl = MUX_s_1_2_2(mux_666_nl, nand_251_nl, or_960_cse);
  assign nand_250_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_85_psp);
  assign mux_668_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_85_psp),
      or_941_cse);
  assign mux_669_nl = MUX_s_1_2_2(nand_250_nl, mux_668_nl, nor_307_cse);
  assign mux_670_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_84_psp),
      or_941_cse);
  assign nand_249_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_84_psp);
  assign mux_671_nl = MUX_s_1_2_2(mux_670_nl, nand_249_nl, or_967_cse);
  assign mux_672_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_83_psp),
      or_941_cse);
  assign nand_248_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_83_psp);
  assign mux_673_nl = MUX_s_1_2_2(mux_672_nl, nand_248_nl, or_967_cse);
  assign nand_247_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_82_psp);
  assign mux_674_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_82_psp),
      or_941_cse);
  assign mux_675_nl = MUX_s_1_2_2(nand_247_nl, mux_674_nl, nor_307_cse);
  assign mux_676_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_81_psp),
      or_941_cse);
  assign nand_246_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_81_psp);
  assign mux_677_nl = MUX_s_1_2_2(mux_676_nl, nand_246_nl, or_960_cse);
  assign nand_245_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_80_psp);
  assign mux_678_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_80_psp),
      or_941_cse);
  assign mux_679_nl = MUX_s_1_2_2(nand_245_nl, mux_678_nl, nor_304_cse);
  assign nand_244_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_79_psp);
  assign mux_680_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_79_psp),
      or_941_cse);
  assign mux_681_nl = MUX_s_1_2_2(nand_244_nl, mux_680_nl, nor_302_cse);
  assign mux_682_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_78_psp),
      or_941_cse);
  assign nand_243_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_78_psp);
  assign mux_683_nl = MUX_s_1_2_2(mux_682_nl, nand_243_nl, or_950_cse);
  assign nand_242_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_77_psp);
  assign mux_684_nl = MUX_s_1_2_2(or_dcpl_56, (~ LOAD_LOOP_for_if_for_for_and_77_psp),
      or_941_cse);
  assign mux_685_nl = MUX_s_1_2_2(nand_242_nl, mux_684_nl, and_3220_cse);
  assign mux_686_nl = MUX_s_1_2_2(or_dcpl_85, (~ LOAD_LOOP_for_if_for_for_and_76_psp),
      or_941_cse);
  assign nand_241_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_76_psp);
  assign mux_687_nl = MUX_s_1_2_2(mux_686_nl, nand_241_nl, or_939_cse);
  assign mux_688_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_75_psp),
      or_941_cse);
  assign nand_333_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_75_psp);
  assign mux_689_nl = MUX_s_1_2_2(mux_688_nl, nand_333_nl, or_939_cse);
  assign nand_332_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_74_psp);
  assign mux_690_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_74_psp),
      or_941_cse);
  assign mux_691_nl = MUX_s_1_2_2(nand_332_nl, mux_690_nl, and_3220_cse);
  assign mux_692_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_73_psp),
      or_941_cse);
  assign nand_240_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_73_psp);
  assign mux_693_nl = MUX_s_1_2_2(mux_692_nl, nand_240_nl, or_950_cse);
  assign nand_239_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_72_psp);
  assign mux_694_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_72_psp),
      or_941_cse);
  assign mux_695_nl = MUX_s_1_2_2(nand_239_nl, mux_694_nl, nor_302_cse);
  assign nand_238_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_71_psp);
  assign mux_696_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_71_psp),
      or_941_cse);
  assign mux_697_nl = MUX_s_1_2_2(nand_238_nl, mux_696_nl, nor_304_cse);
  assign mux_698_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_70_psp),
      or_941_cse);
  assign nand_237_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_70_psp);
  assign mux_699_nl = MUX_s_1_2_2(mux_698_nl, nand_237_nl, or_960_cse);
  assign nand_236_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_69_psp);
  assign mux_700_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_69_psp),
      or_941_cse);
  assign mux_701_nl = MUX_s_1_2_2(nand_236_nl, mux_700_nl, nor_307_cse);
  assign mux_702_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_68_psp),
      or_941_cse);
  assign nand_235_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_68_psp);
  assign mux_703_nl = MUX_s_1_2_2(mux_702_nl, nand_235_nl, or_967_cse);
  assign mux_704_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_67_psp),
      or_941_cse);
  assign nand_234_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_67_psp);
  assign mux_705_nl = MUX_s_1_2_2(mux_704_nl, nand_234_nl, or_967_cse);
  assign nand_233_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_66_psp);
  assign mux_706_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_66_psp),
      or_941_cse);
  assign mux_707_nl = MUX_s_1_2_2(nand_233_nl, mux_706_nl, nor_307_cse);
  assign mux_708_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_65_psp),
      or_941_cse);
  assign nand_232_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_65_psp);
  assign mux_709_nl = MUX_s_1_2_2(mux_708_nl, nand_232_nl, or_960_cse);
  assign nand_231_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_64_psp);
  assign mux_710_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_64_psp),
      or_941_cse);
  assign mux_711_nl = MUX_s_1_2_2(nand_231_nl, mux_710_nl, nor_304_cse);
  assign nand_230_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_63_psp);
  assign mux_712_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_63_psp),
      or_941_cse);
  assign mux_713_nl = MUX_s_1_2_2(nand_230_nl, mux_712_nl, nor_302_cse);
  assign mux_714_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_62_psp),
      or_941_cse);
  assign nand_229_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_62_psp);
  assign mux_715_nl = MUX_s_1_2_2(mux_714_nl, nand_229_nl, or_950_cse);
  assign nand_228_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_61_psp);
  assign mux_716_nl = MUX_s_1_2_2(or_dcpl_66, (~ LOAD_LOOP_for_if_for_for_and_61_psp),
      or_941_cse);
  assign mux_717_nl = MUX_s_1_2_2(nand_228_nl, mux_716_nl, and_3220_cse);
  assign mux_718_nl = MUX_s_1_2_2(or_dcpl_76, (~ LOAD_LOOP_for_if_for_for_and_60_psp),
      or_941_cse);
  assign nand_227_nl = ~(or_941_cse & LOAD_LOOP_for_if_for_for_and_60_psp);
  assign mux_719_nl = MUX_s_1_2_2(mux_718_nl, nand_227_nl, or_939_cse);
  assign and_944_nl = or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 & or_tmp_4;
  assign mux_720_nl = MUX_s_1_2_2(and_tmp_58, and_944_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_943_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_249_psp & or_tmp_4;
  assign mux_721_nl = MUX_s_1_2_2(mux_720_nl, and_943_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_722_nl = MUX_s_1_2_2(mux_721_nl, and_tmp_58, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_694_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_723_nl = MUX_s_1_2_2(and_tmp_61, nor_694_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_946_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_248_psp & or_tmp_4;
  assign mux_724_nl = MUX_s_1_2_2(mux_723_nl, and_946_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_725_nl = MUX_s_1_2_2(mux_724_nl, and_tmp_61, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign and_950_nl = or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 & or_tmp_4;
  assign mux_726_nl = MUX_s_1_2_2(and_tmp_64, and_950_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_949_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_247_psp & or_tmp_4;
  assign mux_727_nl = MUX_s_1_2_2(mux_726_nl, and_949_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_728_nl = MUX_s_1_2_2(mux_727_nl, and_tmp_64, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_693_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_729_nl = MUX_s_1_2_2(and_tmp_67, nor_693_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_952_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_246_psp & or_tmp_4;
  assign mux_730_nl = MUX_s_1_2_2(mux_729_nl, and_952_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_731_nl = MUX_s_1_2_2(mux_730_nl, and_tmp_67, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_692_nl = ~(nand_222_cse | nand_223_cse);
  assign mux_732_nl = MUX_s_1_2_2(and_tmp_70, nor_692_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_955_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_245_psp & or_tmp_4;
  assign mux_733_nl = MUX_s_1_2_2(mux_732_nl, and_955_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_734_nl = MUX_s_1_2_2(mux_733_nl, and_tmp_70, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_691_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_735_nl = MUX_s_1_2_2(and_tmp_73, nor_691_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_958_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_244_psp & or_tmp_4;
  assign mux_736_nl = MUX_s_1_2_2(mux_735_nl, and_958_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_737_nl = MUX_s_1_2_2(mux_736_nl, and_tmp_73, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign and_3209_nl = or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]))
      & or_tmp_4;
  assign mux_738_nl = MUX_s_1_2_2(and_tmp_75, and_3209_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_960_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_243_psp & or_tmp_4;
  assign mux_739_nl = MUX_s_1_2_2(mux_738_nl, and_960_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_740_nl = MUX_s_1_2_2(mux_739_nl, and_tmp_75, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_690_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_741_nl = MUX_s_1_2_2(and_tmp_77, nor_690_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_962_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_242_psp & or_tmp_4;
  assign mux_742_nl = MUX_s_1_2_2(mux_741_nl, and_962_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_743_nl = MUX_s_1_2_2(mux_742_nl, and_tmp_77, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_689_nl = ~(nand_222_cse | nand_224_cse);
  assign mux_744_nl = MUX_s_1_2_2(and_tmp_80, nor_689_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_965_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_241_psp & or_tmp_4;
  assign mux_745_nl = MUX_s_1_2_2(mux_744_nl, and_965_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_746_nl = MUX_s_1_2_2(mux_745_nl, and_tmp_80, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_688_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_218_cse);
  assign mux_747_nl = MUX_s_1_2_2(and_tmp_83, nor_688_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_968_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_240_psp & or_tmp_4;
  assign mux_748_nl = MUX_s_1_2_2(mux_747_nl, and_968_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_749_nl = MUX_s_1_2_2(mux_748_nl, and_tmp_83, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_687_nl = ~(nand_222_cse | nand_225_cse);
  assign mux_750_nl = MUX_s_1_2_2(and_tmp_86, nor_687_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_971_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_239_psp & or_tmp_4;
  assign mux_751_nl = MUX_s_1_2_2(mux_750_nl, and_971_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_752_nl = MUX_s_1_2_2(mux_751_nl, and_tmp_86, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_686_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_215_cse);
  assign mux_753_nl = MUX_s_1_2_2(and_tmp_89, nor_686_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_974_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_238_psp & or_tmp_4;
  assign mux_754_nl = MUX_s_1_2_2(mux_753_nl, and_974_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_755_nl = MUX_s_1_2_2(mux_754_nl, and_tmp_89, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_685_nl = ~(nand_213_cse | nand_214_cse);
  assign mux_756_nl = MUX_s_1_2_2(and_tmp_92, nor_685_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_977_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_237_psp & or_tmp_4;
  assign mux_757_nl = MUX_s_1_2_2(mux_756_nl, and_977_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_758_nl = MUX_s_1_2_2(mux_757_nl, and_tmp_92, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_684_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_212_cse);
  assign mux_759_nl = MUX_s_1_2_2(and_tmp_95, nor_684_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_980_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_236_psp & or_tmp_4;
  assign mux_760_nl = MUX_s_1_2_2(mux_759_nl, and_980_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_761_nl = MUX_s_1_2_2(mux_760_nl, and_tmp_95, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_683_nl = ~(nand_213_cse | nand_212_cse);
  assign mux_762_nl = MUX_s_1_2_2(and_tmp_98, nor_683_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_983_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_235_psp & or_tmp_4;
  assign mux_763_nl = MUX_s_1_2_2(mux_762_nl, and_983_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_764_nl = MUX_s_1_2_2(mux_763_nl, and_tmp_98, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_682_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_214_cse);
  assign mux_765_nl = MUX_s_1_2_2(and_tmp_101, nor_682_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_986_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_234_psp & or_tmp_4;
  assign mux_766_nl = MUX_s_1_2_2(mux_765_nl, and_986_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_767_nl = MUX_s_1_2_2(mux_766_nl, and_tmp_101, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_681_nl = ~(nand_213_cse | nand_215_cse);
  assign mux_768_nl = MUX_s_1_2_2(and_tmp_104, nor_681_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_989_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_233_psp & or_tmp_4;
  assign mux_769_nl = MUX_s_1_2_2(mux_768_nl, and_989_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_770_nl = MUX_s_1_2_2(mux_769_nl, and_tmp_104, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_680_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_225_cse);
  assign mux_771_nl = MUX_s_1_2_2(and_tmp_107, nor_680_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_992_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_232_psp & or_tmp_4;
  assign mux_772_nl = MUX_s_1_2_2(mux_771_nl, and_992_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_773_nl = MUX_s_1_2_2(mux_772_nl, and_tmp_107, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_679_nl = ~(nand_213_cse | nand_218_cse);
  assign mux_774_nl = MUX_s_1_2_2(and_tmp_110, nor_679_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_995_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_231_psp & or_tmp_4;
  assign mux_775_nl = MUX_s_1_2_2(mux_774_nl, and_995_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_776_nl = MUX_s_1_2_2(mux_775_nl, and_tmp_110, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_678_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_224_cse);
  assign mux_777_nl = MUX_s_1_2_2(and_tmp_113, nor_678_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_998_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_230_psp & or_tmp_4;
  assign mux_778_nl = MUX_s_1_2_2(mux_777_nl, and_998_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_779_nl = MUX_s_1_2_2(mux_778_nl, and_tmp_113, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_677_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b111)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_780_nl = MUX_s_1_2_2(and_tmp_116, nor_677_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1001_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_229_psp & or_tmp_4;
  assign mux_781_nl = MUX_s_1_2_2(mux_780_nl, and_1001_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_782_nl = MUX_s_1_2_2(mux_781_nl, and_tmp_116, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_676_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]))
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_783_nl = MUX_s_1_2_2(and_tmp_119, nor_676_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1004_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_228_psp & or_tmp_4;
  assign mux_784_nl = MUX_s_1_2_2(mux_783_nl, and_1004_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_785_nl = MUX_s_1_2_2(mux_784_nl, and_tmp_119, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign and_3208_nl = or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b111)
      & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]))
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]))
      & or_tmp_4;
  assign mux_786_nl = MUX_s_1_2_2(and_tmp_121, and_3208_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1006_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_227_psp & or_tmp_4;
  assign mux_787_nl = MUX_s_1_2_2(mux_786_nl, and_1006_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_788_nl = MUX_s_1_2_2(mux_787_nl, and_tmp_121, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_675_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_223_cse);
  assign mux_789_nl = MUX_s_1_2_2(and_tmp_123, nor_675_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1008_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_226_psp & or_tmp_4;
  assign mux_790_nl = MUX_s_1_2_2(mux_789_nl, and_1008_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_791_nl = MUX_s_1_2_2(mux_790_nl, and_tmp_123, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_674_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b111)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_792_nl = MUX_s_1_2_2(and_tmp_126, nor_674_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1011_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_225_psp & or_tmp_4;
  assign mux_793_nl = MUX_s_1_2_2(mux_792_nl, and_1011_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_794_nl = MUX_s_1_2_2(mux_793_nl, and_tmp_126, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_673_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | nand_199_cse);
  assign mux_795_nl = MUX_s_1_2_2(and_tmp_129, nor_673_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1014_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_224_psp & or_tmp_4;
  assign mux_796_nl = MUX_s_1_2_2(mux_795_nl, and_1014_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_797_nl = MUX_s_1_2_2(mux_796_nl, and_tmp_129, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_672_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b111)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_798_nl = MUX_s_1_2_2(and_tmp_132, nor_672_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1017_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_223_psp & or_tmp_4;
  assign mux_799_nl = MUX_s_1_2_2(mux_798_nl, and_1017_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_800_nl = MUX_s_1_2_2(mux_799_nl, and_tmp_132, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_671_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | nand_197_cse);
  assign mux_801_nl = MUX_s_1_2_2(and_tmp_135, nor_671_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1020_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_222_psp & or_tmp_4;
  assign mux_802_nl = MUX_s_1_2_2(mux_801_nl, and_1020_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_803_nl = MUX_s_1_2_2(mux_802_nl, and_tmp_135, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_670_nl = ~(nand_195_cse | nand_196_cse);
  assign mux_804_nl = MUX_s_1_2_2(and_tmp_138, nor_670_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1023_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_221_psp & or_tmp_4;
  assign mux_805_nl = MUX_s_1_2_2(mux_804_nl, and_1023_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_806_nl = MUX_s_1_2_2(mux_805_nl, and_tmp_138, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_669_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | nand_194_cse);
  assign mux_807_nl = MUX_s_1_2_2(and_tmp_141, nor_669_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1026_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_220_psp & or_tmp_4;
  assign mux_808_nl = MUX_s_1_2_2(mux_807_nl, and_1026_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_809_nl = MUX_s_1_2_2(mux_808_nl, and_tmp_141, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_668_nl = ~(nand_195_cse | nand_194_cse);
  assign mux_810_nl = MUX_s_1_2_2(and_tmp_144, nor_668_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1029_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_219_psp & or_tmp_4;
  assign mux_811_nl = MUX_s_1_2_2(mux_810_nl, and_1029_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_812_nl = MUX_s_1_2_2(mux_811_nl, and_tmp_144, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_667_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b000)
      | nand_196_cse);
  assign mux_813_nl = MUX_s_1_2_2(and_tmp_147, nor_667_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1032_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_218_psp & or_tmp_4;
  assign mux_814_nl = MUX_s_1_2_2(mux_813_nl, and_1032_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_815_nl = MUX_s_1_2_2(mux_814_nl, and_tmp_147, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_666_nl = ~(nand_195_cse | nand_197_cse);
  assign mux_816_nl = MUX_s_1_2_2(and_tmp_150, nor_666_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1035_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_217_psp & or_tmp_4;
  assign mux_817_nl = MUX_s_1_2_2(mux_816_nl, and_1035_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_818_nl = MUX_s_1_2_2(mux_817_nl, and_tmp_150, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_665_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_819_nl = MUX_s_1_2_2(and_tmp_153, nor_665_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1038_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_216_psp & or_tmp_4;
  assign mux_820_nl = MUX_s_1_2_2(mux_819_nl, and_1038_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_821_nl = MUX_s_1_2_2(mux_820_nl, and_tmp_153, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_664_nl = ~(nand_195_cse | nand_199_cse);
  assign mux_822_nl = MUX_s_1_2_2(and_tmp_156, nor_664_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1041_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_215_psp & or_tmp_4;
  assign mux_823_nl = MUX_s_1_2_2(mux_822_nl, and_1041_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_824_nl = MUX_s_1_2_2(mux_823_nl, and_tmp_156, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_663_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_825_nl = MUX_s_1_2_2(and_tmp_159, nor_663_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1044_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_214_psp & or_tmp_4;
  assign mux_826_nl = MUX_s_1_2_2(mux_825_nl, and_1044_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_827_nl = MUX_s_1_2_2(mux_826_nl, and_tmp_159, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_662_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_223_cse);
  assign mux_828_nl = MUX_s_1_2_2(and_tmp_162, nor_662_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1047_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_213_psp & or_tmp_4;
  assign mux_829_nl = MUX_s_1_2_2(mux_828_nl, and_1047_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, and_tmp_162, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_661_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_831_nl = MUX_s_1_2_2(and_tmp_165, nor_661_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1050_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_212_psp & or_tmp_4;
  assign mux_832_nl = MUX_s_1_2_2(mux_831_nl, and_1050_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_833_nl = MUX_s_1_2_2(mux_832_nl, and_tmp_165, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign and_3207_nl = or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b110)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]))
      & or_tmp_4;
  assign mux_834_nl = MUX_s_1_2_2(and_tmp_167, and_3207_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1052_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_211_psp & or_tmp_4;
  assign mux_835_nl = MUX_s_1_2_2(mux_834_nl, and_1052_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_836_nl = MUX_s_1_2_2(mux_835_nl, and_tmp_167, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_660_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_837_nl = MUX_s_1_2_2(and_tmp_169, nor_660_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1054_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_210_psp & or_tmp_4;
  assign mux_838_nl = MUX_s_1_2_2(mux_837_nl, and_1054_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_839_nl = MUX_s_1_2_2(mux_838_nl, and_tmp_169, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_659_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_224_cse);
  assign mux_840_nl = MUX_s_1_2_2(and_tmp_172, nor_659_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1057_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_209_psp & or_tmp_4;
  assign mux_841_nl = MUX_s_1_2_2(mux_840_nl, and_1057_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_842_nl = MUX_s_1_2_2(mux_841_nl, and_tmp_172, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_658_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_218_cse);
  assign mux_843_nl = MUX_s_1_2_2(and_tmp_175, nor_658_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1060_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_208_psp & or_tmp_4;
  assign mux_844_nl = MUX_s_1_2_2(mux_843_nl, and_1060_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_845_nl = MUX_s_1_2_2(mux_844_nl, and_tmp_175, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_657_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_225_cse);
  assign mux_846_nl = MUX_s_1_2_2(and_tmp_178, nor_657_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1063_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_207_psp & or_tmp_4;
  assign mux_847_nl = MUX_s_1_2_2(mux_846_nl, and_1063_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_848_nl = MUX_s_1_2_2(mux_847_nl, and_tmp_178, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_656_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_215_cse);
  assign mux_849_nl = MUX_s_1_2_2(and_tmp_181, nor_656_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1066_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_206_psp & or_tmp_4;
  assign mux_850_nl = MUX_s_1_2_2(mux_849_nl, and_1066_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_851_nl = MUX_s_1_2_2(mux_850_nl, and_tmp_181, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_655_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_214_cse);
  assign mux_852_nl = MUX_s_1_2_2(and_tmp_184, nor_655_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1069_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_205_psp & or_tmp_4;
  assign mux_853_nl = MUX_s_1_2_2(mux_852_nl, and_1069_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_854_nl = MUX_s_1_2_2(mux_853_nl, and_tmp_184, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_654_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_212_cse);
  assign mux_855_nl = MUX_s_1_2_2(and_tmp_187, nor_654_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1072_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_204_psp & or_tmp_4;
  assign mux_856_nl = MUX_s_1_2_2(mux_855_nl, and_1072_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_857_nl = MUX_s_1_2_2(mux_856_nl, and_tmp_187, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_653_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_212_cse);
  assign mux_858_nl = MUX_s_1_2_2(and_tmp_190, nor_653_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1075_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_203_psp & or_tmp_4;
  assign mux_859_nl = MUX_s_1_2_2(mux_858_nl, and_1075_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_860_nl = MUX_s_1_2_2(mux_859_nl, and_tmp_190, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_652_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_214_cse);
  assign mux_861_nl = MUX_s_1_2_2(and_tmp_193, nor_652_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1078_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_202_psp & or_tmp_4;
  assign mux_862_nl = MUX_s_1_2_2(mux_861_nl, and_1078_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_863_nl = MUX_s_1_2_2(mux_862_nl, and_tmp_193, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_651_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_215_cse);
  assign mux_864_nl = MUX_s_1_2_2(and_tmp_196, nor_651_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1081_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_201_psp & or_tmp_4;
  assign mux_865_nl = MUX_s_1_2_2(mux_864_nl, and_1081_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_866_nl = MUX_s_1_2_2(mux_865_nl, and_tmp_196, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_650_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_225_cse);
  assign mux_867_nl = MUX_s_1_2_2(and_tmp_199, nor_650_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1084_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_200_psp & or_tmp_4;
  assign mux_868_nl = MUX_s_1_2_2(mux_867_nl, and_1084_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_869_nl = MUX_s_1_2_2(mux_868_nl, and_tmp_199, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_649_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_218_cse);
  assign mux_870_nl = MUX_s_1_2_2(and_tmp_202, nor_649_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1087_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_199_psp & or_tmp_4;
  assign mux_871_nl = MUX_s_1_2_2(mux_870_nl, and_1087_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_872_nl = MUX_s_1_2_2(mux_871_nl, and_tmp_202, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_648_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_224_cse);
  assign mux_873_nl = MUX_s_1_2_2(and_tmp_205, nor_648_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1090_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_198_psp & or_tmp_4;
  assign mux_874_nl = MUX_s_1_2_2(mux_873_nl, and_1090_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_875_nl = MUX_s_1_2_2(mux_874_nl, and_tmp_205, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_647_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_876_nl = MUX_s_1_2_2(and_tmp_208, nor_647_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1093_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_197_psp & or_tmp_4;
  assign mux_877_nl = MUX_s_1_2_2(mux_876_nl, and_1093_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_878_nl = MUX_s_1_2_2(mux_877_nl, and_tmp_208, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_646_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]))
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_879_nl = MUX_s_1_2_2(and_tmp_211, nor_646_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1096_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_196_psp & or_tmp_4;
  assign mux_880_nl = MUX_s_1_2_2(mux_879_nl, and_1096_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_881_nl = MUX_s_1_2_2(mux_880_nl, and_tmp_211, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_645_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_882_nl = MUX_s_1_2_2(and_tmp_213, nor_645_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1098_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_195_psp & or_tmp_4;
  assign mux_883_nl = MUX_s_1_2_2(mux_882_nl, and_1098_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_884_nl = MUX_s_1_2_2(mux_883_nl, and_tmp_213, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_644_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b001)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_223_cse);
  assign mux_885_nl = MUX_s_1_2_2(and_tmp_215, nor_644_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1100_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_194_psp & or_tmp_4;
  assign mux_886_nl = MUX_s_1_2_2(mux_885_nl, and_1100_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_887_nl = MUX_s_1_2_2(mux_886_nl, and_tmp_215, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_643_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_888_nl = MUX_s_1_2_2(and_tmp_218, nor_643_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1103_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_193_psp & or_tmp_4;
  assign mux_889_nl = MUX_s_1_2_2(mux_888_nl, and_1103_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_890_nl = MUX_s_1_2_2(mux_889_nl, and_tmp_218, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_642_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b00)
      | nand_167_cse);
  assign mux_891_nl = MUX_s_1_2_2(and_tmp_221, nor_642_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1106_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_192_psp & or_tmp_4;
  assign mux_892_nl = MUX_s_1_2_2(mux_891_nl, and_1106_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_893_nl = MUX_s_1_2_2(mux_892_nl, and_tmp_221, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_641_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b110)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_894_nl = MUX_s_1_2_2(and_tmp_224, nor_641_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1109_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_191_psp & or_tmp_4;
  assign mux_895_nl = MUX_s_1_2_2(mux_894_nl, and_1109_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_896_nl = MUX_s_1_2_2(mux_895_nl, and_tmp_224, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_640_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b00)
      | nand_165_cse);
  assign mux_897_nl = MUX_s_1_2_2(and_tmp_227, nor_640_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1112_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_190_psp & or_tmp_4;
  assign mux_898_nl = MUX_s_1_2_2(mux_897_nl, and_1112_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_899_nl = MUX_s_1_2_2(mux_898_nl, and_tmp_227, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_639_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b10)
      | nand_164_cse);
  assign mux_900_nl = MUX_s_1_2_2(and_tmp_230, nor_639_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1115_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_189_psp & or_tmp_4;
  assign mux_901_nl = MUX_s_1_2_2(mux_900_nl, and_1115_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_902_nl = MUX_s_1_2_2(mux_901_nl, and_tmp_230, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_638_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b00)
      | nand_163_cse);
  assign mux_903_nl = MUX_s_1_2_2(and_tmp_233, nor_638_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1118_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_188_psp & or_tmp_4;
  assign mux_904_nl = MUX_s_1_2_2(mux_903_nl, and_1118_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_905_nl = MUX_s_1_2_2(mux_904_nl, and_tmp_233, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_637_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b10)
      | nand_163_cse);
  assign mux_906_nl = MUX_s_1_2_2(and_tmp_236, nor_637_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1121_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_187_psp & or_tmp_4;
  assign mux_907_nl = MUX_s_1_2_2(mux_906_nl, and_1121_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_908_nl = MUX_s_1_2_2(mux_907_nl, and_tmp_236, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_636_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b00)
      | nand_164_cse);
  assign mux_909_nl = MUX_s_1_2_2(and_tmp_239, nor_636_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1124_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_186_psp & or_tmp_4;
  assign mux_910_nl = MUX_s_1_2_2(mux_909_nl, and_1124_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_911_nl = MUX_s_1_2_2(mux_910_nl, and_tmp_239, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_635_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b10)
      | nand_165_cse);
  assign mux_912_nl = MUX_s_1_2_2(and_tmp_242, nor_635_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1127_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_185_psp & or_tmp_4;
  assign mux_913_nl = MUX_s_1_2_2(mux_912_nl, and_1127_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_914_nl = MUX_s_1_2_2(mux_913_nl, and_tmp_242, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_634_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_915_nl = MUX_s_1_2_2(and_tmp_245, nor_634_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1130_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_184_psp & or_tmp_4;
  assign mux_916_nl = MUX_s_1_2_2(mux_915_nl, and_1130_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_917_nl = MUX_s_1_2_2(mux_916_nl, and_tmp_245, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_633_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2:1]!=2'b10)
      | nand_167_cse);
  assign mux_918_nl = MUX_s_1_2_2(and_tmp_248, nor_633_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1133_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_183_psp & or_tmp_4;
  assign mux_919_nl = MUX_s_1_2_2(mux_918_nl, and_1133_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_920_nl = MUX_s_1_2_2(mux_919_nl, and_tmp_248, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_632_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_921_nl = MUX_s_1_2_2(and_tmp_251, nor_632_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1136_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_182_psp & or_tmp_4;
  assign mux_922_nl = MUX_s_1_2_2(mux_921_nl, and_1136_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_923_nl = MUX_s_1_2_2(mux_922_nl, and_tmp_251, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_631_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_223_cse);
  assign mux_924_nl = MUX_s_1_2_2(and_tmp_254, nor_631_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1139_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_181_psp & or_tmp_4;
  assign mux_925_nl = MUX_s_1_2_2(mux_924_nl, and_1139_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_926_nl = MUX_s_1_2_2(mux_925_nl, and_tmp_254, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_630_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_927_nl = MUX_s_1_2_2(and_tmp_257, nor_630_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1142_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_180_psp & or_tmp_4;
  assign mux_928_nl = MUX_s_1_2_2(mux_927_nl, and_1142_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_929_nl = MUX_s_1_2_2(mux_928_nl, and_tmp_257, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign and_3206_nl = or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b101)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]))
      & or_tmp_4;
  assign mux_930_nl = MUX_s_1_2_2(and_tmp_259, and_3206_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1144_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_179_psp & or_tmp_4;
  assign mux_931_nl = MUX_s_1_2_2(mux_930_nl, and_1144_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_932_nl = MUX_s_1_2_2(mux_931_nl, and_tmp_259, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_629_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_933_nl = MUX_s_1_2_2(and_tmp_261, nor_629_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1146_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_178_psp & or_tmp_4;
  assign mux_934_nl = MUX_s_1_2_2(mux_933_nl, and_1146_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_935_nl = MUX_s_1_2_2(mux_934_nl, and_tmp_261, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_628_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_224_cse);
  assign mux_936_nl = MUX_s_1_2_2(and_tmp_264, nor_628_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1149_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_177_psp & or_tmp_4;
  assign mux_937_nl = MUX_s_1_2_2(mux_936_nl, and_1149_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_938_nl = MUX_s_1_2_2(mux_937_nl, and_tmp_264, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_627_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_218_cse);
  assign mux_939_nl = MUX_s_1_2_2(and_tmp_267, nor_627_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1152_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_176_psp & or_tmp_4;
  assign mux_940_nl = MUX_s_1_2_2(mux_939_nl, and_1152_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_941_nl = MUX_s_1_2_2(mux_940_nl, and_tmp_267, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_626_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_225_cse);
  assign mux_942_nl = MUX_s_1_2_2(and_tmp_270, nor_626_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1155_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_175_psp & or_tmp_4;
  assign mux_943_nl = MUX_s_1_2_2(mux_942_nl, and_1155_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_944_nl = MUX_s_1_2_2(mux_943_nl, and_tmp_270, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_625_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_215_cse);
  assign mux_945_nl = MUX_s_1_2_2(and_tmp_273, nor_625_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1158_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_174_psp & or_tmp_4;
  assign mux_946_nl = MUX_s_1_2_2(mux_945_nl, and_1158_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_947_nl = MUX_s_1_2_2(mux_946_nl, and_tmp_273, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_624_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_214_cse);
  assign mux_948_nl = MUX_s_1_2_2(and_tmp_276, nor_624_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1161_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_173_psp & or_tmp_4;
  assign mux_949_nl = MUX_s_1_2_2(mux_948_nl, and_1161_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_950_nl = MUX_s_1_2_2(mux_949_nl, and_tmp_276, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_623_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_212_cse);
  assign mux_951_nl = MUX_s_1_2_2(and_tmp_279, nor_623_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1164_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_172_psp & or_tmp_4;
  assign mux_952_nl = MUX_s_1_2_2(mux_951_nl, and_1164_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_953_nl = MUX_s_1_2_2(mux_952_nl, and_tmp_279, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_622_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_212_cse);
  assign mux_954_nl = MUX_s_1_2_2(and_tmp_282, nor_622_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1167_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_171_psp & or_tmp_4;
  assign mux_955_nl = MUX_s_1_2_2(mux_954_nl, and_1167_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_956_nl = MUX_s_1_2_2(mux_955_nl, and_tmp_282, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_621_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_214_cse);
  assign mux_957_nl = MUX_s_1_2_2(and_tmp_285, nor_621_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1170_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_170_psp & or_tmp_4;
  assign mux_958_nl = MUX_s_1_2_2(mux_957_nl, and_1170_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_959_nl = MUX_s_1_2_2(mux_958_nl, and_tmp_285, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_620_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_215_cse);
  assign mux_960_nl = MUX_s_1_2_2(and_tmp_288, nor_620_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1173_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_169_psp & or_tmp_4;
  assign mux_961_nl = MUX_s_1_2_2(mux_960_nl, and_1173_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_962_nl = MUX_s_1_2_2(mux_961_nl, and_tmp_288, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_619_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_225_cse);
  assign mux_963_nl = MUX_s_1_2_2(and_tmp_291, nor_619_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1176_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_168_psp & or_tmp_4;
  assign mux_964_nl = MUX_s_1_2_2(mux_963_nl, and_1176_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_965_nl = MUX_s_1_2_2(mux_964_nl, and_tmp_291, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_618_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_218_cse);
  assign mux_966_nl = MUX_s_1_2_2(and_tmp_294, nor_618_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1179_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_167_psp & or_tmp_4;
  assign mux_967_nl = MUX_s_1_2_2(mux_966_nl, and_1179_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_968_nl = MUX_s_1_2_2(mux_967_nl, and_tmp_294, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_617_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_224_cse);
  assign mux_969_nl = MUX_s_1_2_2(and_tmp_297, nor_617_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1182_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_166_psp & or_tmp_4;
  assign mux_970_nl = MUX_s_1_2_2(mux_969_nl, and_1182_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_971_nl = MUX_s_1_2_2(mux_970_nl, and_tmp_297, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_616_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_972_nl = MUX_s_1_2_2(and_tmp_300, nor_616_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1185_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_165_psp & or_tmp_4;
  assign mux_973_nl = MUX_s_1_2_2(mux_972_nl, and_1185_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_974_nl = MUX_s_1_2_2(mux_973_nl, and_tmp_300, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_615_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]))
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_975_nl = MUX_s_1_2_2(and_tmp_303, nor_615_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1188_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_164_psp & or_tmp_4;
  assign mux_976_nl = MUX_s_1_2_2(mux_975_nl, and_1188_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_977_nl = MUX_s_1_2_2(mux_976_nl, and_tmp_303, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_614_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_978_nl = MUX_s_1_2_2(and_tmp_305, nor_614_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1190_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_163_psp & or_tmp_4;
  assign mux_979_nl = MUX_s_1_2_2(mux_978_nl, and_1190_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_980_nl = MUX_s_1_2_2(mux_979_nl, and_tmp_305, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_613_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_223_cse);
  assign mux_981_nl = MUX_s_1_2_2(and_tmp_307, nor_613_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1192_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_162_psp & or_tmp_4;
  assign mux_982_nl = MUX_s_1_2_2(mux_981_nl, and_1192_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_983_nl = MUX_s_1_2_2(mux_982_nl, and_tmp_307, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_612_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_984_nl = MUX_s_1_2_2(and_tmp_310, nor_612_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1195_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_161_psp & or_tmp_4;
  assign mux_985_nl = MUX_s_1_2_2(mux_984_nl, and_1195_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_986_nl = MUX_s_1_2_2(mux_985_nl, and_tmp_310, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_611_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | nand_199_cse);
  assign mux_987_nl = MUX_s_1_2_2(and_tmp_313, nor_611_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1198_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_160_psp & or_tmp_4;
  assign mux_988_nl = MUX_s_1_2_2(mux_987_nl, and_1198_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_989_nl = MUX_s_1_2_2(mux_988_nl, and_tmp_313, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_610_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b101)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_990_nl = MUX_s_1_2_2(and_tmp_316, nor_610_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1201_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_159_psp & or_tmp_4;
  assign mux_991_nl = MUX_s_1_2_2(mux_990_nl, and_1201_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_992_nl = MUX_s_1_2_2(mux_991_nl, and_tmp_316, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_609_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | nand_197_cse);
  assign mux_993_nl = MUX_s_1_2_2(and_tmp_319, nor_609_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1204_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_158_psp & or_tmp_4;
  assign mux_994_nl = MUX_s_1_2_2(mux_993_nl, and_1204_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_995_nl = MUX_s_1_2_2(mux_994_nl, and_tmp_319, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_608_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | nand_196_cse);
  assign mux_996_nl = MUX_s_1_2_2(and_tmp_322, nor_608_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1207_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_157_psp & or_tmp_4;
  assign mux_997_nl = MUX_s_1_2_2(mux_996_nl, and_1207_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_998_nl = MUX_s_1_2_2(mux_997_nl, and_tmp_322, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_607_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | nand_194_cse);
  assign mux_999_nl = MUX_s_1_2_2(and_tmp_325, nor_607_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1210_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_156_psp & or_tmp_4;
  assign mux_1000_nl = MUX_s_1_2_2(mux_999_nl, and_1210_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1001_nl = MUX_s_1_2_2(mux_1000_nl, and_tmp_325, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_606_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | nand_194_cse);
  assign mux_1002_nl = MUX_s_1_2_2(and_tmp_328, nor_606_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1213_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_155_psp & or_tmp_4;
  assign mux_1003_nl = MUX_s_1_2_2(mux_1002_nl, and_1213_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1004_nl = MUX_s_1_2_2(mux_1003_nl, and_tmp_328, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_605_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b010)
      | nand_196_cse);
  assign mux_1005_nl = MUX_s_1_2_2(and_tmp_331, nor_605_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1216_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_154_psp & or_tmp_4;
  assign mux_1006_nl = MUX_s_1_2_2(mux_1005_nl, and_1216_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1007_nl = MUX_s_1_2_2(mux_1006_nl, and_tmp_331, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_604_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | nand_197_cse);
  assign mux_1008_nl = MUX_s_1_2_2(and_tmp_334, nor_604_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1219_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_153_psp & or_tmp_4;
  assign mux_1009_nl = MUX_s_1_2_2(mux_1008_nl, and_1219_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1010_nl = MUX_s_1_2_2(mux_1009_nl, and_tmp_334, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_603_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_1011_nl = MUX_s_1_2_2(and_tmp_337, nor_603_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1222_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_152_psp & or_tmp_4;
  assign mux_1012_nl = MUX_s_1_2_2(mux_1011_nl, and_1222_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1013_nl = MUX_s_1_2_2(mux_1012_nl, and_tmp_337, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_602_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | nand_199_cse);
  assign mux_1014_nl = MUX_s_1_2_2(and_tmp_340, nor_602_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1225_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_151_psp & or_tmp_4;
  assign mux_1015_nl = MUX_s_1_2_2(mux_1014_nl, and_1225_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1016_nl = MUX_s_1_2_2(mux_1015_nl, and_tmp_340, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_601_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_1017_nl = MUX_s_1_2_2(and_tmp_343, nor_601_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1228_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_150_psp & or_tmp_4;
  assign mux_1018_nl = MUX_s_1_2_2(mux_1017_nl, and_1228_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1019_nl = MUX_s_1_2_2(mux_1018_nl, and_tmp_343, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_600_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_223_cse);
  assign mux_1020_nl = MUX_s_1_2_2(and_tmp_346, nor_600_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1231_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_149_psp & or_tmp_4;
  assign mux_1021_nl = MUX_s_1_2_2(mux_1020_nl, and_1231_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1022_nl = MUX_s_1_2_2(mux_1021_nl, and_tmp_346, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_599_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_1023_nl = MUX_s_1_2_2(and_tmp_349, nor_599_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1234_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_148_psp & or_tmp_4;
  assign mux_1024_nl = MUX_s_1_2_2(mux_1023_nl, and_1234_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1025_nl = MUX_s_1_2_2(mux_1024_nl, and_tmp_349, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_598_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1]))
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_1026_nl = MUX_s_1_2_2(and_tmp_351, nor_598_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1236_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_147_psp & or_tmp_4;
  assign mux_1027_nl = MUX_s_1_2_2(mux_1026_nl, and_1236_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1028_nl = MUX_s_1_2_2(mux_1027_nl, and_tmp_351, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_597_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_1029_nl = MUX_s_1_2_2(and_tmp_353, nor_597_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1238_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_146_psp & or_tmp_4;
  assign mux_1030_nl = MUX_s_1_2_2(mux_1029_nl, and_1238_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1031_nl = MUX_s_1_2_2(mux_1030_nl, and_tmp_353, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_596_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_224_cse);
  assign mux_1032_nl = MUX_s_1_2_2(and_tmp_356, nor_596_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1241_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_145_psp & or_tmp_4;
  assign mux_1033_nl = MUX_s_1_2_2(mux_1032_nl, and_1241_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1034_nl = MUX_s_1_2_2(mux_1033_nl, and_tmp_356, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_595_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_218_cse);
  assign mux_1035_nl = MUX_s_1_2_2(and_tmp_359, nor_595_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1244_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_144_psp & or_tmp_4;
  assign mux_1036_nl = MUX_s_1_2_2(mux_1035_nl, and_1244_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1037_nl = MUX_s_1_2_2(mux_1036_nl, and_tmp_359, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_594_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_225_cse);
  assign mux_1038_nl = MUX_s_1_2_2(and_tmp_362, nor_594_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1247_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_143_psp & or_tmp_4;
  assign mux_1039_nl = MUX_s_1_2_2(mux_1038_nl, and_1247_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1040_nl = MUX_s_1_2_2(mux_1039_nl, and_tmp_362, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_593_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_215_cse);
  assign mux_1041_nl = MUX_s_1_2_2(and_tmp_365, nor_593_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1250_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_142_psp & or_tmp_4;
  assign mux_1042_nl = MUX_s_1_2_2(mux_1041_nl, and_1250_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1043_nl = MUX_s_1_2_2(mux_1042_nl, and_tmp_365, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_592_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_214_cse);
  assign mux_1044_nl = MUX_s_1_2_2(and_tmp_368, nor_592_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1253_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_141_psp & or_tmp_4;
  assign mux_1045_nl = MUX_s_1_2_2(mux_1044_nl, and_1253_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1046_nl = MUX_s_1_2_2(mux_1045_nl, and_tmp_368, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_591_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_212_cse);
  assign mux_1047_nl = MUX_s_1_2_2(and_tmp_371, nor_591_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1256_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_140_psp & or_tmp_4;
  assign mux_1048_nl = MUX_s_1_2_2(mux_1047_nl, and_1256_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1049_nl = MUX_s_1_2_2(mux_1048_nl, and_tmp_371, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_590_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_212_cse);
  assign mux_1050_nl = MUX_s_1_2_2(and_tmp_374, nor_590_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1259_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_139_psp & or_tmp_4;
  assign mux_1051_nl = MUX_s_1_2_2(mux_1050_nl, and_1259_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1052_nl = MUX_s_1_2_2(mux_1051_nl, and_tmp_374, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_589_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_214_cse);
  assign mux_1053_nl = MUX_s_1_2_2(and_tmp_377, nor_589_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1262_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_138_psp & or_tmp_4;
  assign mux_1054_nl = MUX_s_1_2_2(mux_1053_nl, and_1262_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1055_nl = MUX_s_1_2_2(mux_1054_nl, and_tmp_377, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_588_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_215_cse);
  assign mux_1056_nl = MUX_s_1_2_2(and_tmp_380, nor_588_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1265_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_137_psp & or_tmp_4;
  assign mux_1057_nl = MUX_s_1_2_2(mux_1056_nl, and_1265_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1058_nl = MUX_s_1_2_2(mux_1057_nl, and_tmp_380, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_587_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_225_cse);
  assign mux_1059_nl = MUX_s_1_2_2(and_tmp_383, nor_587_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1268_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_136_psp & or_tmp_4;
  assign mux_1060_nl = MUX_s_1_2_2(mux_1059_nl, and_1268_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1061_nl = MUX_s_1_2_2(mux_1060_nl, and_tmp_383, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_586_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | nand_218_cse);
  assign mux_1062_nl = MUX_s_1_2_2(and_tmp_386, nor_586_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1271_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_135_psp & or_tmp_4;
  assign mux_1063_nl = MUX_s_1_2_2(mux_1062_nl, and_1271_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1064_nl = MUX_s_1_2_2(mux_1063_nl, and_tmp_386, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_585_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_224_cse);
  assign mux_1065_nl = MUX_s_1_2_2(and_tmp_389, nor_585_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1274_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_134_psp & or_tmp_4;
  assign mux_1066_nl = MUX_s_1_2_2(mux_1065_nl, and_1274_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1067_nl = MUX_s_1_2_2(mux_1066_nl, and_tmp_389, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_584_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_223_cse);
  assign mux_1068_nl = MUX_s_1_2_2(and_tmp_392, nor_584_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1277_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_133_psp & or_tmp_4;
  assign mux_1069_nl = MUX_s_1_2_2(mux_1068_nl, and_1277_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1070_nl = MUX_s_1_2_2(mux_1069_nl, and_tmp_392, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign and_3205_nl = or_9_cse & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3==3'b011)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (~ (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0]))
      & or_tmp_4;
  assign mux_1071_nl = MUX_s_1_2_2(and_tmp_395, and_3205_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1280_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_132_psp & or_tmp_4;
  assign mux_1072_nl = MUX_s_1_2_2(mux_1071_nl, and_1280_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1073_nl = MUX_s_1_2_2(mux_1072_nl, and_tmp_395, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_583_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      | (~ LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      | (~ or_tmp_4));
  assign mux_1074_nl = MUX_s_1_2_2(and_tmp_397, nor_583_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1282_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_131_psp & or_tmp_4;
  assign mux_1075_nl = MUX_s_1_2_2(mux_1074_nl, and_1282_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1076_nl = MUX_s_1_2_2(mux_1075_nl, and_tmp_397, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_582_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b011)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b10)
      | nand_223_cse);
  assign mux_1077_nl = MUX_s_1_2_2(and_tmp_399, nor_582_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1284_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_130_psp & or_tmp_4;
  assign mux_1078_nl = MUX_s_1_2_2(mux_1077_nl, and_1284_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1079_nl = MUX_s_1_2_2(mux_1078_nl, and_tmp_399, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_581_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_224_cse);
  assign mux_1080_nl = MUX_s_1_2_2(and_tmp_402, nor_581_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1287_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_129_psp & or_tmp_4;
  assign mux_1081_nl = MUX_s_1_2_2(mux_1080_nl, and_1287_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1082_nl = MUX_s_1_2_2(mux_1081_nl, and_tmp_402, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_580_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      | (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_0_sva_1 & or_tmp_4)));
  assign mux_1083_nl = MUX_s_1_2_2(and_tmp_405, nor_580_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1290_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_128_psp & or_tmp_4;
  assign mux_1084_nl = MUX_s_1_2_2(mux_1083_nl, and_1290_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1085_nl = MUX_s_1_2_2(mux_1084_nl, and_tmp_405, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_579_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3!=3'b100)
      | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1!=2'b00)
      | nand_225_cse);
  assign mux_1086_nl = MUX_s_1_2_2(and_tmp_408, nor_579_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1293_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_127_psp & or_tmp_4;
  assign mux_1087_nl = MUX_s_1_2_2(mux_1086_nl, and_1293_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1088_nl = MUX_s_1_2_2(mux_1087_nl, and_tmp_408, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_578_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      | (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_1_sva_1 & or_tmp_4)));
  assign mux_1089_nl = MUX_s_1_2_2(and_tmp_411, nor_578_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1296_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_126_psp & or_tmp_4;
  assign mux_1090_nl = MUX_s_1_2_2(mux_1089_nl, and_1296_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1091_nl = MUX_s_1_2_2(mux_1090_nl, and_tmp_411, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_577_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      | (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1==2'b11)
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_3_sva_1 & or_tmp_4)));
  assign mux_1092_nl = MUX_s_1_2_2(and_tmp_414, nor_577_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1299_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_125_psp & or_tmp_4;
  assign mux_1093_nl = MUX_s_1_2_2(mux_1092_nl, and_1299_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1094_nl = MUX_s_1_2_2(mux_1093_nl, and_tmp_414, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign nor_576_nl = ~((~ or_9_cse) | (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[2])
      | (~((LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_5_3[1:0]==2'b11)
      & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[1])
      & LOAD_LOOP_for_if_2_for_for_and_stg_1_2_sva_1 & (LOAD_LOOP_for_if_2_for_for_LOAD_LOOP_for_if_2_for_for_conc_decb_6_1_sva_2_2_1[0])
      & or_tmp_4)));
  assign mux_1095_nl = MUX_s_1_2_2(and_tmp_417, nor_576_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_2);
  assign and_1302_nl = or_tmp_853 & LOAD_LOOP_for_if_2_for_for_and_124_psp & or_tmp_4;
  assign mux_1096_nl = MUX_s_1_2_2(mux_1095_nl, and_1302_nl, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[1]);
  assign mux_1097_nl = MUX_s_1_2_2(mux_1096_nl, and_tmp_417, lfst_exit_LOAD_LOOP_for_if_2_for_lpi_2_dfm_st_2_1_0[0]);
  assign LOAD_LOOP_for_if_2_for_for_if_index_in_mux_8_nl = MUX_v_8_2_2(({3'b000 ,
      LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1}), (conf_info_rsci_idat_mxwt[103:96]),
      fsm_output[1]);
  assign LOAD_LOOP_for_if_2_for_for_if_index_in_mux_9_nl = MUX_v_8_2_2(({n_w_in_acc_psp_sva
      , (conf_info_crt_sva_231_0[192])}), (conf_info_rsci_idat_mxwt[103:96]), fsm_output[1]);
  assign z_out_15_0 = conv_u2u_16_16(LOAD_LOOP_for_if_2_for_for_if_index_in_mux_8_nl
      * LOAD_LOOP_for_if_2_for_for_if_index_in_mux_9_nl);
  assign LOAD_LOOP_for_if_2_for_for_if_index_in_mux_10_nl = MUX_v_8_2_2(({n_h_in_acc_psp_sva
      , (conf_info_crt_sva_231_0[160])}), (conf_info_rsci_idat_mxwt[39:32]), fsm_output[1]);
  assign operator_43_true_and_1_nl = (z_out_10[16]) & (z_out_10[0]);
  assign nl_operator_43_true_operator_43_true_acc_1_nl = (z_out_10[8:1]) + conv_u2s_1_8(operator_43_true_and_1_nl);
  assign operator_43_true_operator_43_true_acc_1_nl = nl_operator_43_true_operator_43_true_acc_1_nl[7:0];
  assign LOAD_LOOP_for_if_2_for_for_if_index_in_mux_11_nl = MUX_v_13_2_2((z_out_15_0[12:0]),
      (signext_13_8(operator_43_true_operator_43_true_acc_1_nl)), fsm_output[1]);
  assign nl_z_out_1 = LOAD_LOOP_for_if_2_for_for_if_index_in_mux_10_nl * LOAD_LOOP_for_if_2_for_for_if_index_in_mux_11_nl;
  assign z_out_1 = nl_z_out_1[13:0];
  assign batch_size_mux1h_14_nl = MUX1HOT_v_8_3_2((conf_info_rsci_idat_mxwt[135:128]),
      ({3'b000 , LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1}), (conf_info_crt_sva_231_0[199:192]),
      {(fsm_output[1]) , and_3316_cse , and_3318_cse});
  assign batch_size_mux1h_15_nl = MUX1HOT_v_16_3_2(z_out_15_0, batch_size_mul_4_cse_sva,
      ({11'b00000000000 , LOAD_LOOP_for_k_5_0_lpi_2_dfm_4_0_1}), {(fsm_output[1])
      , and_3316_cse , and_3318_cse});
  assign nl_z_out_2_15_0 = batch_size_mux1h_14_nl * batch_size_mux1h_15_nl;
  assign z_out_2_15_0 = nl_z_out_2_15_0[15:0];
  assign LOAD_LOOP_for_if_for_for_index_f_mux_2_nl = MUX_v_8_2_2(({5'b00000 , LOAD_LOOP_for_if_for_m_2_0_lpi_2_mx1}),
      (conf_info_rsci_idat_mxwt[199:192]), fsm_output[1]);
  assign LOAD_LOOP_for_if_for_for_index_f_mux_3_nl = MUX_v_8_2_2(({2'b00 , (conf_info_crt_sva_231_0[101:96])}),
      (conf_info_rsci_idat_mxwt[167:160]), fsm_output[1]);
  assign z_out_3_15_0 = conv_u2u_16_16(LOAD_LOOP_for_if_for_for_index_f_mux_2_nl
      * LOAD_LOOP_for_if_for_for_index_f_mux_3_nl);
  assign pad_mux_5_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[7:0]), (conf_info_crt_sva_231_0[167:160]),
      fsm_output[2]);
  assign pad_mux_6_nl = MUX_v_14_2_2(({{5{z_out_13[8]}}, z_out_13}), ({1'b0 , (z_out_2_15_0[12:0])}),
      fsm_output[2]);
  assign nl_z_out_4 = $signed(conv_u2s_8_9(pad_mux_5_nl)) * $signed(pad_mux_6_nl);
  assign z_out_4 = nl_z_out_4[16:0];
  assign LOAD_LOOP_for_mux_13_nl = MUX_v_8_2_2(({3'b000 , LOAD_LOOP_fl_5_0_sva_4_0}),
      (conf_info_rsci_idat_mxwt[71:64]), fsm_output[1]);
  assign LOAD_LOOP_for_mux_14_nl = MUX_v_16_2_2(batch_size_mul_3_cse_sva, z_out_2_15_0,
      fsm_output[1]);
  assign nl_z_out_5 = LOAD_LOOP_for_mux_13_nl * LOAD_LOOP_for_mux_14_nl;
  assign z_out_5 = nl_z_out_5[15:0];
  assign batch_size_mux_7_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[135:128]), ({4'b0000
      , LOAD_BATCH_LOOP_b_4_0_sva_3_0}), fsm_output[2]);
  assign batch_size_mux_8_nl = MUX_v_16_2_2(z_out_3_15_0, batch_size_sva, fsm_output[2]);
  assign nl_z_out_6 = batch_size_mux_7_nl * batch_size_mux_8_nl;
  assign z_out_6 = nl_z_out_6[15:0];
  assign operator_8_false_1_mux_4_nl = MUX_v_2_2_2(({1'b1 , (z_out_8[0])}), (z_out_9[1:0]),
      and_3338_cse);
  assign operator_8_false_1_operator_8_false_1_nor_1_nl = ~((z_out_8[2]) | and_3338_cse);
  assign operator_8_false_1_mux_5_nl = MUX_s_1_2_2((~ (z_out_8[1])), (z_out_9[2]),
      and_3338_cse);
  assign nl_acc_nl = conv_u2u_3_4({operator_8_false_1_mux_4_nl , operator_8_false_1_operator_8_false_1_nor_1_nl})
      + conv_u2u_2_4({operator_8_false_1_mux_5_nl , 1'b1});
  assign acc_nl = nl_acc_nl[3:0];
  assign z_out_7 = readslicef_4_3_1(acc_nl);
  assign operator_8_false_1_mux_6_nl = MUX_v_2_2_2(({1'b0 , (operator_8_false_1_acc_psp_sva_1[0])}),
      (~ (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[3:2])), and_3338_cse);
  assign operator_8_false_1_mux_7_nl = MUX_v_2_2_2((~ (operator_8_false_1_acc_psp_sva_1[2:1])),
      ({1'b0 , (LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[4])}), and_3338_cse);
  assign nl_acc_1_nl = conv_u2u_3_4({operator_8_false_1_mux_6_nl , 1'b1}) + conv_s2u_3_4({operator_8_false_1_mux_7_nl
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[3:0];
  assign z_out_8 = readslicef_4_3_1(acc_1_nl);
  assign nl_operator_8_false_3_acc_4_nl = ({(~ (operator_8_false_3_acc_psp_sva_1[2]))
      , 2'b00}) + conv_s2u_1_3(operator_8_false_3_acc_psp_sva_1[3]) + conv_u2u_1_3(operator_8_false_3_acc_psp_sva_1[2]);
  assign operator_8_false_3_acc_4_nl = nl_operator_8_false_3_acc_4_nl[2:0];
  assign operator_8_false_2_mux_3_nl = MUX_v_3_2_2(z_out_8, operator_8_false_3_acc_4_nl,
      or_tmp_2431);
  assign operator_8_false_2_mux_4_nl = MUX_v_2_2_2((LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1[1:0]),
      (operator_8_false_3_acc_psp_sva_1[1:0]), or_tmp_2431);
  assign nl_z_out_9 = operator_8_false_2_mux_3_nl + ({1'b1 , operator_8_false_2_mux_4_nl});
  assign z_out_9 = nl_z_out_9[2:0];
  assign LOAD_LOOP_for_LOAD_LOOP_for_and_2_nl = (z_out_4[16]) & (~(and_3316_cse |
      and_3318_cse));
  assign LOAD_LOOP_for_LOAD_LOOP_for_mux_5_nl = MUX_v_16_2_2(z_out_12, (z_out_4[15:0]),
      fsm_output[1]);
  assign LOAD_LOOP_for_mux1h_9_nl = MUX1HOT_v_16_3_2(z_out_6, ({{7{z_out_11[8]}},
      z_out_11}), LOAD_LOOP_for_mul_cse_lpi_2, {and_3316_cse , (fsm_output[1]) ,
      and_3318_cse});
  assign nl_z_out_10 = ({LOAD_LOOP_for_LOAD_LOOP_for_and_2_nl , LOAD_LOOP_for_LOAD_LOOP_for_mux_5_nl})
      + conv_s2u_16_17(LOAD_LOOP_for_mux1h_9_nl);
  assign z_out_10 = nl_z_out_10[16:0];
  assign pad_pad_pad_nor_1_nl = ~(MUX_v_3_2_2((conf_info_rsci_idat_mxwt[199:197]),
      3'b111, (fsm_output[2])));
  assign pad_mux_7_nl = MUX_v_5_2_2((~ (conf_info_rsci_idat_mxwt[196:192])), LOAD_LOOP_for_if_2_for_row_4_0_lpi_2_mx1,
      fsm_output[2]);
  assign pad_mux_8_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[103:96]), (~ pad_sva),
      fsm_output[2]);
  assign nl_acc_4_nl = ({1'b1 , pad_pad_pad_nor_1_nl , pad_mux_7_nl , 1'b1}) + conv_u2u_9_10({pad_mux_8_nl
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[9:0];
  assign z_out_11 = readslicef_10_9_1(acc_4_nl);
  assign batch_size_mux1h_16_nl = MUX1HOT_v_16_3_2(z_out_6, z_out_5, batch_size_mul_2_cse_sva,
      {(fsm_output[1]) , and_3316_cse , and_3318_cse});
  assign batch_size_mux1h_17_nl = MUX1HOT_v_16_3_2(z_out_5, z_out_2_15_0, (z_out_4[15:0]),
      {(fsm_output[1]) , and_3316_cse , and_3318_cse});
  assign nl_z_out_12 = batch_size_mux1h_16_nl + batch_size_mux1h_17_nl;
  assign z_out_12 = nl_z_out_12[15:0];
  assign operator_8_false_3_mux_1_nl = MUX_v_8_2_2((conf_info_crt_sva_231_0[103:96]),
      (conf_info_rsci_idat_mxwt[199:192]), fsm_output[1]);
  assign nl_z_out_13 = conv_u2u_8_9(operator_8_false_3_mux_1_nl) + 9'b111111111;
  assign z_out_13 = nl_z_out_13[8:0];

  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input [0:0] sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] readslicef_10_9_1;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_10_9_1 = tmp[8:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [2:0] readslicef_4_3_1;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_4_3_1 = tmp[2:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [12:0] signext_13_8;
    input [7:0] vector;
  begin
    signext_13_8= {{5{vector[7]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input [0:0] vector;
  begin
    signext_5_1= {{4{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] conv_s2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_3 = {vector[1], vector};
  end
  endfunction


  function automatic [3:0] conv_s2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [2:0] conv_s2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_3 = {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_s2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2u_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [9:0] conv_s2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [2:0] conv_u2s_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_3 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_3_6 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_6 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_5_8 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_8 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_5_13 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_13 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_13_13 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_13 = vector;
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_16 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute_core
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, buf_linear_rsc_dat,
      buf_linear_rsc_vld, buf_linear_rsc_rdy, plm_kernel_rsc_dat, plm_kernel_rsc_vld,
      plm_kernel_rsc_rdy, var_output_rsc_dat, var_output_rsc_vld, var_output_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input [4031:0] buf_linear_rsc_dat;
  input buf_linear_rsc_vld;
  output buf_linear_rsc_rdy;
  input [1567:0] plm_kernel_rsc_dat;
  input plm_kernel_rsc_vld;
  output plm_kernel_rsc_rdy;
  output [31:0] var_output_rsc_dat;
  output var_output_rsc_vld;
  input var_output_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire core_wen;
  wire conf_info_rsci_bawt;
  wire conf_info_rsci_wen_comp;
  wire [63:0] conf_info_rsci_idat_mxwt;
  wire buf_linear_rsci_bawt;
  wire buf_linear_rsci_wen_comp;
  wire [4031:0] buf_linear_rsci_idat_mxwt;
  wire plm_kernel_rsci_bawt;
  wire plm_kernel_rsci_wen_comp;
  wire [1567:0] plm_kernel_rsci_idat_mxwt;
  wire var_output_rsci_bawt;
  wire var_output_rsci_wen_comp;
  wire done_rsci_bawt;
  wire done_rsci_wen_comp;
  reg var_output_rsci_idat_31;
  reg [29:0] var_output_rsci_idat_30_1;
  reg var_output_rsci_idat_0;
  wire [4:0] COMPUTE_LOOP_acc_tmp;
  wire [5:0] nl_COMPUTE_LOOP_acc_tmp;
  wire [8:0] operator_8_false_8_acc_tmp;
  wire [9:0] nl_operator_8_false_8_acc_tmp;
  wire [5:0] CONVOLUTION_LOOP_acc_tmp;
  wire [6:0] nl_CONVOLUTION_LOOP_acc_tmp;
  wire [8:0] operator_8_false_7_acc_tmp;
  wire [9:0] nl_operator_8_false_7_acc_tmp;
  wire [5:0] CONVOLUTION_LOOP_for_acc_tmp;
  wire [6:0] nl_CONVOLUTION_LOOP_for_acc_tmp;
  wire CONVOLUTION_LOOP_for_if_equal_tmp;
  wire CONVOLUTION_LOOP_for_for_if_CONVOLUTION_LOOP_for_for_if_nand_tmp;
  wire [8:0] operator_8_false_5_acc_tmp;
  wire [9:0] nl_operator_8_false_5_acc_tmp;
  wire [8:0] operator_8_false_4_acc_tmp;
  wire [9:0] nl_operator_8_false_4_acc_tmp;
  wire [8:0] operator_8_false_3_acc_tmp;
  wire [9:0] nl_operator_8_false_3_acc_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp;
  wire [8:0] operator_8_false_1_acc_tmp;
  wire [9:0] nl_operator_8_false_1_acc_tmp;
  wire or_dcpl_11;
  wire or_dcpl_12;
  wire and_dcpl_8;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire mux_tmp_27;
  wire mux_tmp_28;
  wire and_dcpl_25;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_tmp_13;
  wire mux_tmp_29;
  wire and_dcpl_34;
  wire or_dcpl_32;
  wire or_dcpl_33;
  wire or_dcpl_36;
  wire or_dcpl_38;
  wire or_dcpl_42;
  wire and_tmp_14;
  wire not_tmp_46;
  wire and_dcpl_40;
  wire and_tmp_28;
  wire nand_tmp_20;
  wire and_tmp_29;
  wire and_dcpl_47;
  wire or_dcpl_51;
  wire and_dcpl_54;
  wire or_dcpl_57;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire or_dcpl_62;
  wire or_dcpl_63;
  wire not_tmp_91;
  wire or_dcpl_64;
  wire or_dcpl_75;
  wire or_dcpl_76;
  wire and_dcpl_61;
  wire and_dcpl_66;
  wire and_dcpl_68;
  wire and_dcpl_71;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0;
  wire lfst_exit_CONVOLUTION_LOOP_1_lpi_1_dfm_1;
  wire exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0;
  wire exitL_exit_COMPUTE_LOOP_sva_mx0;
  wire exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0;
  reg [3:0] COMPUTE_LOOP_b_4_0_lpi_1_dfm_1_3_0;
  wire exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0w0;
  wire exit_CONVOLUTION_LOOP_sva_3;
  reg [4:0] CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_1_4_0;
  wire exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_2_mx0w0;
  wire exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0;
  reg [4:0] CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_4;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1;
  wire CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_56_1;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1_dfm_1_mx0;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_64_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_65_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_66_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_6_67_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_5_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_67_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_66_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_65_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_64_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_stg_7_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1;
  reg [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1;
  reg COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1;
  wire CONVOLUTION_LOOP_for_for_for_acc_56_sva_2;
  wire [54:0] CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2;
  wire CONVOLUTION_LOOP_for_for_for_acc_0_sva_2;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1;
  reg [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_1_dfm_1;
  wire [57:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_5_psp_sva_1;
  wire [58:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_5_psp_sva_1;
  wire [63:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_1_sdt_sva_1;
  wire unequal_tmp_1;
  reg exitL_exit_COMPUTE_LOOP_sva;
  wire exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1;
  reg main_stage_v_1;
  reg exit_COMPUTE_LOOP_lpi_1_dfm_3_st_2;
  reg main_stage_v_3;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1;
  reg main_stage_v_2;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1;
  reg COMPUTE_LOOP_asn_itm_1;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1;
  reg exit_COMPUTE_LOOP_lpi_1_dfm_3_st_1;
  wire exit_COMPUTE_LOOP_lpi_1_dfm_3_mx0w0;
  reg exit_COMPUTE_LOOP_lpi_1_dfm_1;
  reg exit_CONVOLUTION_LOOP_lpi_1_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_sva_2_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_sva_2;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2;
  wire [54:0] CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_55_1_1;
  wire [57:0] CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1;
  wire [58:0] nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1;
  wire [57:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1;
  wire [58:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1;
  reg reg_done_rsci_iswt0_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_6_cse;
  reg reg_var_output_rsci_iswt0_cse;
  reg reg_conf_info_rsci_iswt0_cse;
  reg reg_plm_kernel_rsci_iswt0_cse;
  reg reg_buf_linear_rsci_iswt0_cse;
  wire COMPUTE_LOOP_and_2_cse;
  wire COMPUTE_LOOP_buf_tmp_acc_data_and_cse;
  wire or_41_cse;
  wire nand_74_cse;
  wire and_156_cse;
  wire or_59_cse;
  wire or_57_cse;
  wire or_58_cse;
  wire nand_76_cse;
  wire or_61_cse;
  wire asn_done_rsci_oswt_and_cse;
  wire and_6_cse;
  wire nor_42_cse;
  wire nor_32_cse;
  wire or_289_cse;
  wire or_290_cse;
  wire nand_52_cse;
  wire or_155_cse;
  wire or_157_cse;
  wire or_163_cse;
  wire mux_50_cse;
  wire exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
  wire [4:0] CONVOLUTION_LOOP_for_for_i_4_0_sva_2;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2;
  wire [3:0] nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_1;
  wire [2:0] z_out;
  wire [1:0] z_out_1;
  wire [7:0] z_out_5;
  wire [8:0] nl_z_out_5;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_1;
  reg [6:0] CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1;
  reg [7:0] n_w_out_lpi_1_dfm_1;
  reg [7:0] n_h_out_lpi_1_dfm_1;
  reg [1567:0] COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm;
  reg [4031:0] COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm;
  reg [6:0] CONVOLUTION_LOOP_for_for_for_y_mul_cse_6_0_lpi_1_dfm;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_1;
  reg CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1;
  reg [54:0] CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1;
  reg [7:0] conf_info_crt_lpi_1_dfm_231_224;
  reg [7:0] conf_info_crt_lpi_1_dfm_135_128;
  reg [7:0] conf_info_crt_lpi_1_dfm_103_96;
  reg [7:0] conf_info_crt_lpi_1_dfm_71_64;
  reg [7:0] conf_info_crt_lpi_1_dfm_7_0;
  wire [7:0] if_acc_4_cse_1;
  wire [8:0] nl_if_acc_4_cse_1;
  wire [7:0] pad_sva_1;
  wire signed [16:0] nl_pad_sva_1;
  wire [10:0] else_acc_2_psp_sva_1;
  wire [11:0] nl_else_acc_2_psp_sva_1;
  wire [9:0] else_acc_4_cse_1;
  wire [10:0] nl_else_acc_4_cse_1;
  wire [10:0] else_acc_psp_sva_1;
  wire [11:0] nl_else_acc_psp_sva_1;
  wire [16:0] pad_acc_psp_sva_1;
  wire [17:0] nl_pad_acc_psp_sva_1;
  wire [7:0] conf_info_crt_lpi_1_dfm_7_0_mx0;
  wire [1:0] operator_8_false_1_acc_imod_2_sva_1;
  wire [3:0] nl_operator_8_false_1_acc_imod_2_sva_1;
  wire [2:0] operator_8_false_1_acc_imod_1_sva_1;
  wire [3:0] nl_operator_8_false_1_acc_imod_1_sva_1;
  wire [3:0] operator_8_false_1_acc_imod_sva_1;
  wire [4:0] nl_operator_8_false_1_acc_imod_sva_1;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_for_asn_2929_mx0w0;
  wire [12:0] nl_CONVOLUTION_LOOP_for_for_for_for_asn_2929_mx0w0;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0;
  wire [2:0] operator_8_false_2_acc_psp_1;
  wire [3:0] nl_operator_8_false_2_acc_psp_1;
  wire [3:0] operator_8_false_2_acc_5_sdt_1;
  wire [5:0] nl_operator_8_false_2_acc_5_sdt_1;
  wire [4:0] operator_8_false_3_acc_imod_sva_1;
  wire [5:0] nl_operator_8_false_3_acc_imod_sva_1;
  wire [7:0] conf_info_crt_lpi_1_dfm_231_224_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_71_64_mx0;
  wire [7:0] n_w_out_lpi_1_dfm_2;
  wire CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1;
  wire [54:0] CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1_dfm_1_mx0;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1_dfm_2;
  wire [54:0] COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1_dfm_2;
  wire [7:0] n_h_out_lpi_1_dfm_2;
  wire [7:0] conf_info_crt_lpi_1_dfm_135_128_mx0;
  wire CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2;
  wire [3:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2;
  wire [7:0] conf_info_crt_lpi_1_dfm_103_96_mx0;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1;
  wire [4031:0] COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_for_x_tmp_2_0_lpi_1_dfm_1;
  wire [6:0] CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0;
  wire [11:0] nl_CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0;
  wire [6:0] CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1_dfm_mx0;
  wire [1567:0] COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0;
  wire COMPUTE_LOOP_asn_itm_1_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_2_rgt;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_3_rgt;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_5_rgt;
  wire COMPUTE_LOOP_or_2_cse;
  wire or_314_cse;
  wire operator_8_false_5_acc_itm_3_1;
  wire operator_8_false_6_acc_itm_3_1;
  wire operator_8_false_3_acc_itm_4_1;
  wire operator_8_false_4_acc_itm_4_1;
  wire mux_66_cse_1;
  wire [2:0] z_out_2_2_0;
  wire [3:0] nl_z_out_2_2_0;

  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl;
  wire[29:0] CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] and_159_nl;
  wire[0:0] and_149_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] or_135_nl;
  wire[0:0] nand_26_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] or_184_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_not_339_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_not_14_nl;
  wire[0:0] COMPUTE_LOOP_not_19_nl;
  wire[4:0] CONVOLUTION_LOOP_CONVOLUTION_LOOP_CONVOLUTION_LOOP_mux_nl;
  wire[0:0] COMPUTE_LOOP_COMPUTE_LOOP_COMPUTE_LOOP_COMPUTE_LOOP_not_1_nl;
  wire[4:0] CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_mux_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_not_22_nl;
  wire[2:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_4_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_not_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_not_26_nl;
  wire[0:0] COMPUTE_LOOP_mux_4_nl;
  wire[0:0] CONVOLUTION_LOOP_mux_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_mux_6_nl;
  wire[7:0] operator_43_true_operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_operator_43_true_acc_nl;
  wire[0:0] operator_43_true_and_nl;
  wire[8:0] pad_acc_2_nl;
  wire[9:0] nl_pad_acc_2_nl;
  wire[16:0] pad_mul_nl;
  wire signed [17:0] nl_pad_mul_nl;
  wire[8:0] operator_8_false_acc_nl;
  wire[9:0] nl_operator_8_false_acc_nl;
  wire[1:0] operator_8_false_1_acc_8_nl;
  wire[2:0] nl_operator_8_false_1_acc_8_nl;
  wire[1:0] operator_8_false_1_acc_7_nl;
  wire[2:0] nl_operator_8_false_1_acc_7_nl;
  wire[2:0] operator_8_false_1_acc_6_nl;
  wire[4:0] nl_operator_8_false_1_acc_6_nl;
  wire[1:0] operator_8_false_1_acc_4_nl;
  wire[3:0] nl_operator_8_false_1_acc_4_nl;
  wire[3:0] operator_8_false_3_acc_4_nl;
  wire[4:0] nl_operator_8_false_3_acc_4_nl;
  wire[8:0] acc_3_nl;
  wire[9:0] nl_acc_3_nl;
  wire[7:0] if_mux_4_nl;
  wire[7:0] if_mux_5_nl;
  wire[0:0] operator_42_true_and_1_nl;
  wire[54:0] CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl;
  wire[54:0] CONVOLUTION_LOOP_for_for_for_else_nor_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_nl;
  wire[54:0] CONVOLUTION_LOOP_for_for_for_else_mux_972_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_973_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_972_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_976_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_973_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_978_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_975_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_976_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_984_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_977_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_978_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_988_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_979_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_981_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_996_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_983_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_984_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_985_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_987_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_988_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_989_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_991_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_993_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_995_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_996_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_997_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_999_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1297_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1626_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1628_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1299_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1630_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1300_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1632_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1301_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1634_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1636_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1303_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1638_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1304_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1640_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1305_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1642_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1306_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1644_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1307_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1646_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1308_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1648_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1309_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1650_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1652_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1311_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1654_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1312_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1656_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1313_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1658_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1660_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1315_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1662_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1316_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1664_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1317_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1666_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1318_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1668_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1319_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1670_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1320_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1672_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1321_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1674_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1676_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1323_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1678_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1324_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1680_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1325_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1682_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1326_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1684_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1327_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1686_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1328_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1688_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1329_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1690_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1330_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1692_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1331_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1694_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1332_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1696_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1333_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1698_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1334_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1700_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1335_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1702_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1336_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1704_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1337_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1706_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1338_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1708_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1339_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1710_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1340_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1712_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1341_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1714_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1342_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1716_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1343_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1718_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1344_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1720_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1345_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1722_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1346_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1724_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1347_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1726_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1348_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1728_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1349_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1730_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1350_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1732_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1351_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1734_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1352_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1736_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1353_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1738_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1354_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1740_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1355_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1742_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1356_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1744_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1357_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1746_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1358_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1748_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1359_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1750_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1360_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1752_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1361_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1754_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1362_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1756_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1363_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1758_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1364_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1760_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1365_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1762_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1366_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1764_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1367_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1766_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1368_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1768_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1369_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1770_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1370_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1772_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1371_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1774_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1372_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1776_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1373_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1778_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1374_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1780_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1375_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1782_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1376_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1784_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1377_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1786_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1378_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1788_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1379_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1790_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1380_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1792_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1381_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1794_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1382_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1796_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1383_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1798_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1384_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1800_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1385_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1802_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1386_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1804_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1387_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1806_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1388_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1808_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1389_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1810_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1390_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1812_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1391_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1814_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1392_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1816_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1393_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1818_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1394_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1820_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1395_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1822_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1396_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1824_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1397_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1826_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1398_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1828_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1399_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1830_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1400_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1832_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1401_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1834_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1402_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1836_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1403_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1838_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1404_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1840_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1405_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1842_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1406_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1844_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1407_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1846_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1408_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1848_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1409_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1850_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1410_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1852_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1411_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1854_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1412_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1856_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1413_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1858_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1414_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1860_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1415_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1862_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1416_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1864_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1417_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1866_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1418_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1868_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1419_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1870_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1420_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1872_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1421_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1874_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1422_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1876_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1423_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1878_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1424_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1880_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1425_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1882_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1426_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1884_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1427_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1886_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1428_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1888_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1429_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1890_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1430_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1892_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1431_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1894_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1432_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1896_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1433_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1898_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1434_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1900_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1435_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1902_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1436_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1904_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1437_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1906_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1438_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1908_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1439_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1910_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1440_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1912_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1441_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1914_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1442_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1916_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1443_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1918_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1444_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1920_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1445_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1922_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1446_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1924_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1447_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1926_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1448_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1928_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1449_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1930_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1450_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1932_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1451_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1934_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1452_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1936_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1453_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1938_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1454_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1940_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1455_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1942_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1456_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1944_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1457_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1946_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1458_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1948_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1459_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1950_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1460_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1952_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1461_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1954_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1462_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1956_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1463_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1958_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1464_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1960_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1465_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1962_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1466_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1964_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1467_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1966_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1468_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1968_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1469_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1970_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1470_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1972_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1471_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1472_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1976_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1473_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1978_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1474_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1475_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1476_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1984_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1477_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1478_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1988_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1479_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1480_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1481_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1482_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1996_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1483_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1484_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2000_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1485_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1486_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1487_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1488_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2008_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1489_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2012_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1491_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1492_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1493_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1494_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2020_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1495_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1496_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2024_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1497_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1498_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1499_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1500_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2032_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1501_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1502_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2036_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1503_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1504_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1505_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1506_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2044_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1507_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1508_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2048_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1509_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1510_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1511_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1512_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2056_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1513_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1514_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2060_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1515_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1516_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1517_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1518_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2068_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1519_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1520_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2072_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1521_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1522_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1523_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1524_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2080_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1525_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1526_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2084_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1527_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1528_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1529_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1530_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2092_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1531_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1532_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2096_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1533_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1534_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1535_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1536_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1537_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1538_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1539_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1540_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1541_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1542_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1543_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1544_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1545_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1546_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1547_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1548_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1549_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1550_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1551_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1552_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1553_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1554_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1555_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1556_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1557_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1558_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1559_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1560_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1561_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1562_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1563_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1564_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1565_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1566_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1567_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1568_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1569_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1570_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1571_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1572_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1573_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1574_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1575_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1576_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1577_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1578_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1579_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1580_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1581_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1582_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1583_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1584_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1585_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1586_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1587_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1588_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1589_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1590_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1591_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1592_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1593_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1594_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1595_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1596_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1597_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1598_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1599_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1600_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1601_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1602_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1603_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1604_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1605_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1606_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1607_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1608_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1609_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1610_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1611_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1612_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1613_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1614_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1615_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1616_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1617_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1618_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_2268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1619_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_2_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_3_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_6_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_7_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_2_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_10_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_11_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_3_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_14_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_15_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_4_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_18_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_19_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_5_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_22_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_23_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_6_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_26_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_27_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_7_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_30_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_31_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_8_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_34_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_35_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_9_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_38_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_39_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_10_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_42_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_43_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_11_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_46_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_47_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_12_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_50_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_51_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_13_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_54_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_55_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_14_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_58_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_59_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_15_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_62_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_63_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_16_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_66_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_67_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_17_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_70_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_71_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_18_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_74_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_75_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_19_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_78_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_79_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_20_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_82_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_83_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_21_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_86_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_87_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_22_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_90_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_91_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_23_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_94_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_95_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_24_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_98_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_99_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_25_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_103_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_26_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_107_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_27_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_111_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_28_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_115_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_29_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_119_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_30_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_123_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_31_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_127_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_32_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_131_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_33_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_135_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_34_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_139_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_35_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_143_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_36_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_147_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_37_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_151_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_38_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_155_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_39_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_159_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_40_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_163_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_41_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_167_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_42_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_171_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_43_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_175_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_44_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_179_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_45_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_183_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_46_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_187_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_47_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_191_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_48_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_195_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_49_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_199_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_50_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_203_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_51_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_207_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_52_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_211_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_53_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_215_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_54_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_219_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_55_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_223_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_56_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_227_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_57_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_231_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_58_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_235_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_59_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_239_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_60_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_243_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_61_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_247_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_62_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_251_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_63_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_255_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_64_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_259_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_65_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_263_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_66_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_267_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_67_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_271_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_68_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_275_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_69_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_279_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_70_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_283_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_71_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_287_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_72_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_291_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_73_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_295_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_74_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_299_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_75_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_303_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_76_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_306_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_307_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_77_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_311_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_78_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_315_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_79_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_318_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_319_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_80_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_323_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_81_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_326_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_327_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_82_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_330_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_331_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_83_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_334_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_335_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_84_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_338_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_339_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_85_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_342_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_343_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_86_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_346_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_347_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_87_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_350_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_351_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_88_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_354_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_355_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_89_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_358_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_359_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_90_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_362_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_363_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_91_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_366_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_367_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_92_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_370_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_371_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_93_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_374_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_375_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_94_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_378_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_379_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_95_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_382_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_383_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_96_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_386_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_387_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_97_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_390_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_391_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_98_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_394_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_395_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_99_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_398_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_399_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_402_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_403_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_101_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_406_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_407_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_410_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_411_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_103_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_414_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_415_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_418_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_419_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_105_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_422_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_423_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_426_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_427_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_107_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_430_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_431_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_434_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_435_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_109_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_438_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_439_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_442_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_443_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_111_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_446_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_447_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_450_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_451_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_113_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_454_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_455_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_458_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_459_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_115_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_462_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_463_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_466_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_467_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_117_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_470_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_471_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_474_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_475_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_119_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_478_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_479_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_482_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_483_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_121_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_486_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_487_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_491_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_123_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_494_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_495_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_498_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_499_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_125_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_502_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_503_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_506_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_507_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_127_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_510_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_511_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_514_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_515_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_129_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_518_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_519_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_522_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_523_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_131_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_526_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_527_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_530_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_531_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_133_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_534_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_535_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_538_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_539_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_135_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_542_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_543_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_546_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_547_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_137_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_550_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_551_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_554_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_555_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_139_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_558_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_559_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_562_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_563_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_141_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_566_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_567_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_570_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_571_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_143_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_574_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_575_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_578_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_579_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_145_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_582_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_583_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_586_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_587_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_147_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_590_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_591_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_594_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_595_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_149_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_598_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_599_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_602_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_603_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_151_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_606_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_607_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_610_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_611_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_153_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_614_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_615_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_618_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_619_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_155_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_622_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_623_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_626_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_627_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_157_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_630_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_631_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_634_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_635_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_159_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_638_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_639_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_642_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_643_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_161_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_646_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_647_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_650_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_651_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_163_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_654_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_655_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_658_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_659_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_165_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_662_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_663_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_666_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_667_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_167_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_670_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_671_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_674_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_675_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_169_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_678_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_679_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_682_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_683_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_171_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_686_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_687_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_690_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_691_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_173_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_694_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_695_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_698_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_699_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_175_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_702_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_703_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_706_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_707_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_177_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_710_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_711_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_714_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_715_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_179_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_718_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_719_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_722_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_723_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_181_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_726_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_727_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_730_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_731_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_183_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_734_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_735_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_738_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_739_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_185_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_742_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_743_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_746_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_747_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_187_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_750_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_751_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_754_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_755_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_189_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_758_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_759_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_762_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_763_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_191_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_766_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_767_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_770_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_771_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_193_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_774_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_775_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_778_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_779_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_195_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_782_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_783_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_786_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_787_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_197_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_790_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_791_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_794_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_795_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_199_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_798_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_799_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_802_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_803_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_201_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_806_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_807_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_810_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_811_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_203_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_814_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_815_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_818_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_819_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_205_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_822_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_823_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_826_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_827_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_207_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_830_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_831_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_834_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_835_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_209_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_838_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_839_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_842_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_843_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_211_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_846_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_847_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_850_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_851_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_213_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_854_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_855_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_858_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_859_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_215_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_862_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_863_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_866_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_867_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_217_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_870_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_871_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_874_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_875_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_219_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_878_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_879_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_882_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_883_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_221_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_886_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_887_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_890_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_891_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_223_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_894_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_895_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_898_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_899_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_225_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_902_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_903_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_906_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_907_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_227_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_910_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_911_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_914_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_915_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_229_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_918_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_919_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_922_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_923_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_231_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_926_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_927_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_930_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_931_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_233_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_934_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_935_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_938_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_939_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_235_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_942_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_943_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_946_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_947_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_237_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_950_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_951_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_954_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_955_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_239_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_958_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_959_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_962_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_963_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_241_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_966_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_967_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_970_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_971_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_243_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_975_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_978_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_979_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_245_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_983_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_987_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_247_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_991_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_995_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_249_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_999_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1003_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_251_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1007_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1011_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_253_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1015_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1019_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_255_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1023_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1027_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_257_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1031_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1035_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_259_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1039_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1043_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_261_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1047_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1051_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_263_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1055_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1059_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_265_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1063_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1067_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_267_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1071_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1075_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_269_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1079_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1083_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_271_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1087_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1091_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_273_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1095_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1099_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_275_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1103_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_276_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1107_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_277_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1111_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1115_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_279_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1119_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1123_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_281_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1127_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1131_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_283_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1135_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1139_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_285_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1143_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1147_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_287_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1151_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_288_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1155_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_289_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1159_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1163_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_291_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1167_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1171_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_293_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1175_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1179_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_295_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1183_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1187_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_297_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1191_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1195_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_299_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1199_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_300_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1203_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_301_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1207_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1211_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_303_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1215_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_304_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1219_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_305_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1223_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_306_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1227_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_307_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1231_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_308_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1235_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_309_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1239_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1243_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_311_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1247_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_312_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1251_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_313_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1255_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1259_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_315_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1263_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_316_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1267_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_317_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1271_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_318_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1275_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_319_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1279_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_320_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1283_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_321_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1287_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1291_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_or_323_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_and_1295_nl;
  wire[8:0] acc_4_nl;
  wire[9:0] nl_acc_4_nl;
  wire[7:0] if_mux_6_nl;
  wire[7:0] if_mux_7_nl;
  wire[0:0] operator_42_true_1_and_1_nl;
  wire[3:0] operator_8_false_5_acc_nl;
  wire[4:0] nl_operator_8_false_5_acc_nl;
  wire[3:0] operator_8_false_6_acc_nl;
  wire[4:0] nl_operator_8_false_6_acc_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_and_nl;
  wire[31:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_7_nl;
  wire[5:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_nl;
  wire[6:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_nl;
  wire[31:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_8_nl;
  wire[5:0] CONVOLUTION_LOOP_for_for_for_for_for_index_f_acc_nl;
  wire[6:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_index_f_acc_nl;
  wire[5:0] CONVOLUTION_LOOP_for_for_for_for_for_index_f_mul_nl;
  wire[8:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_index_f_mul_nl;
  wire[2:0] CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_mux1h_7_nl;
  wire[1:0] operator_8_false_1_acc_3_nl;
  wire[2:0] nl_operator_8_false_1_acc_3_nl;
  wire[2:0] operator_8_false_2_acc_2_nl;
  wire[3:0] nl_operator_8_false_2_acc_2_nl;
  wire[2:0] operator_8_false_3_operator_8_false_3_acc_nl;
  wire[3:0] nl_operator_8_false_3_operator_8_false_3_acc_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_and_3_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_nand_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] and_62_nl;
  wire[0:0] mux_49_nl;
  wire[0:0] and_60_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] and_143_nl;
  wire[0:0] and_144_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] nand_46_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] or_244_nl;
  wire[0:0] nand_47_nl;
  wire[4:0] operator_8_false_3_acc_nl;
  wire[5:0] nl_operator_8_false_3_acc_nl;
  wire[4:0] operator_8_false_4_acc_nl;
  wire[5:0] nl_operator_8_false_4_acc_nl;
  wire[3:0] acc_nl;
  wire[4:0] nl_acc_nl;
  wire[1:0] operator_8_false_2_mux_4_nl;
  wire[0:0] operator_8_false_2_and_1_nl;
  wire[1:0] operator_8_false_2_mux_5_nl;
  wire[2:0] acc_1_nl;
  wire[3:0] nl_acc_1_nl;
  wire[0:0] operator_8_false_1_mux_2_nl;
  wire[0:0] operator_8_false_1_and_1_nl;
  wire[0:0] operator_8_false_1_mux_3_nl;
  wire[2:0] operator_8_false_2_mux_6_nl;
  wire[2:0] operator_8_false_3_acc_7_nl;
  wire[4:0] nl_operator_8_false_3_acc_7_nl;
  wire[2:0] operator_8_false_2_mux_7_nl;
  wire[1:0] operator_8_false_2_acc_7_nl;
  wire[2:0] nl_operator_8_false_2_acc_7_nl;
  wire[7:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_9_nl;
  wire[0:0] nand_85_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_compute_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg;
  assign nl_compute_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg = ~(or_dcpl_42
      | (~(conf_info_rsci_bawt & COMPUTE_LOOP_asn_itm_1)) | and_dcpl_31 | or_dcpl_38);
  wire [0:0] nl_compute_core_buf_linear_rsci_inst_buf_linear_rsci_oswt_unreg;
  assign nl_compute_core_buf_linear_rsci_inst_buf_linear_rsci_oswt_unreg = ~(or_dcpl_42
      | or_dcpl_51 | (~(buf_linear_rsci_bawt & exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1
      & main_stage_v_1)));
  wire [0:0] nl_compute_core_plm_kernel_rsci_inst_plm_kernel_rsci_oswt_unreg;
  assign nl_compute_core_plm_kernel_rsci_inst_plm_kernel_rsci_oswt_unreg = ~(or_dcpl_42
      | and_dcpl_32 | (~(plm_kernel_rsci_bawt & exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1))
      | or_dcpl_38);
  wire [0:0] nl_compute_core_var_output_rsci_inst_var_output_rsci_oswt_unreg;
  assign nl_compute_core_var_output_rsci_inst_var_output_rsci_oswt_unreg = ~(and_6_cse
      | (~ var_output_rsci_bawt) | (~(CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1 & main_stage_v_2)));
  wire [31:0] nl_compute_core_var_output_rsci_inst_var_output_rsci_idat;
  assign nl_compute_core_var_output_rsci_inst_var_output_rsci_idat = {var_output_rsci_idat_31
      , var_output_rsci_idat_30_1 , var_output_rsci_idat_0};
  esp_acc_conv2dlb_cxx_catapult_compute_core_conf_info_rsci compute_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(nl_compute_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg[0:0]),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_iswt0(reg_conf_info_rsci_iswt0_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_buf_linear_rsci compute_core_buf_linear_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .buf_linear_rsc_dat(buf_linear_rsc_dat),
      .buf_linear_rsc_vld(buf_linear_rsc_vld),
      .buf_linear_rsc_rdy(buf_linear_rsc_rdy),
      .core_wen(core_wen),
      .buf_linear_rsci_oswt_unreg(nl_compute_core_buf_linear_rsci_inst_buf_linear_rsci_oswt_unreg[0:0]),
      .buf_linear_rsci_bawt(buf_linear_rsci_bawt),
      .buf_linear_rsci_iswt0(reg_buf_linear_rsci_iswt0_cse),
      .buf_linear_rsci_wen_comp(buf_linear_rsci_wen_comp),
      .buf_linear_rsci_idat_mxwt(buf_linear_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_plm_kernel_rsci compute_core_plm_kernel_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_kernel_rsc_dat(plm_kernel_rsc_dat),
      .plm_kernel_rsc_vld(plm_kernel_rsc_vld),
      .plm_kernel_rsc_rdy(plm_kernel_rsc_rdy),
      .core_wen(core_wen),
      .plm_kernel_rsci_oswt_unreg(nl_compute_core_plm_kernel_rsci_inst_plm_kernel_rsci_oswt_unreg[0:0]),
      .plm_kernel_rsci_bawt(plm_kernel_rsci_bawt),
      .plm_kernel_rsci_iswt0(reg_plm_kernel_rsci_iswt0_cse),
      .plm_kernel_rsci_wen_comp(plm_kernel_rsci_wen_comp),
      .plm_kernel_rsci_idat_mxwt(plm_kernel_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_var_output_rsci compute_core_var_output_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .var_output_rsc_dat(var_output_rsc_dat),
      .var_output_rsc_vld(var_output_rsc_vld),
      .var_output_rsc_rdy(var_output_rsc_rdy),
      .core_wen(core_wen),
      .var_output_rsci_oswt_unreg(nl_compute_core_var_output_rsci_inst_var_output_rsci_oswt_unreg[0:0]),
      .var_output_rsci_bawt(var_output_rsci_bawt),
      .var_output_rsci_iswt0(reg_var_output_rsci_iswt0_cse),
      .var_output_rsci_wen_comp(var_output_rsci_wen_comp),
      .var_output_rsci_idat(nl_compute_core_var_output_rsci_inst_var_output_rsci_idat[31:0])
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_done_rsci compute_core_done_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(asn_done_rsci_oswt_and_cse),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_iswt0(reg_done_rsci_iswt0_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_compute_core_staller compute_core_staller_inst (
      .core_wen(core_wen),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .buf_linear_rsci_wen_comp(buf_linear_rsci_wen_comp),
      .plm_kernel_rsci_wen_comp(plm_kernel_rsci_wen_comp),
      .var_output_rsci_wen_comp(var_output_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  assign asn_done_rsci_oswt_and_cse = done_rsci_bawt & exit_COMPUTE_LOOP_lpi_1_dfm_3_st_2
      & main_stage_v_3;
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_6_cse = core_wen & (~(or_dcpl_36 |
      (~ CONVOLUTION_LOOP_for_if_equal_tmp) | (operator_8_false_3_acc_tmp[8:5]!=4'b0000)
      | or_dcpl_33));
  assign or_155_cse = (~((~((COMPUTE_LOOP_b_4_0_lpi_1_dfm_1_3_0 == (operator_8_false_8_acc_tmp[3:0]))
      & (operator_8_false_8_acc_tmp[7:4]==4'b0000))) | (operator_8_false_8_acc_tmp[8])))
      | (COMPUTE_LOOP_acc_tmp[4]);
  assign or_157_cse = exit_CONVOLUTION_LOOP_sva_3 | (CONVOLUTION_LOOP_acc_tmp[5]);
  assign or_163_cse = nor_32_cse | (CONVOLUTION_LOOP_for_acc_tmp[5]);
  assign nand_52_cse = ~(or_289_cse & operator_8_false_3_acc_itm_4_1);
  assign COMPUTE_LOOP_and_2_cse = core_wen & (~(or_dcpl_42 | and_dcpl_32 | or_dcpl_33));
  assign and_6_cse = (~ done_rsci_bawt) & exit_COMPUTE_LOOP_lpi_1_dfm_3_st_2 & main_stage_v_3;
  assign and_156_cse = core_wen & (~ or_dcpl_57);
  assign COMPUTE_LOOP_buf_tmp_acc_data_and_cse = core_wen & (~(or_dcpl_36 | or_dcpl_33));
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_2_rgt = (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1)
      & and_dcpl_66;
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_3_rgt = exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1
      & and_dcpl_66;
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_5_rgt = exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1
      & and_dcpl_73;
  assign or_41_cse = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)
      | (operator_8_false_1_acc_tmp[8]);
  assign nor_42_cse = ~((~ operator_8_false_6_acc_itm_3_1) | CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp);
  assign or_290_cse = (~((CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1 == (operator_8_false_4_acc_tmp[4:0]))
      & (operator_8_false_4_acc_tmp[7:5]==3'b000))) | (operator_8_false_4_acc_tmp[8]);
  assign nand_74_cse = ~(or_290_cse & operator_8_false_4_acc_itm_4_1);
  assign or_289_cse = CONVOLUTION_LOOP_for_for_if_CONVOLUTION_LOOP_for_for_if_nand_tmp
      | (operator_8_false_5_acc_tmp[8]);
  assign or_59_cse = (~ COMPUTE_LOOP_asn_itm_1) | conf_info_rsci_bawt;
  assign or_57_cse = (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1) |
      buf_linear_rsci_bawt;
  assign or_58_cse = (~ exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1) | plm_kernel_rsci_bawt;
  assign exitL_exit_COMPUTE_LOOP_sva_mx0 = MUX_s_1_2_2(exitL_exit_COMPUTE_LOOP_sva,
      exit_COMPUTE_LOOP_lpi_1_dfm_3_mx0w0, main_stage_v_1);
  assign COMPUTE_LOOP_mux_4_nl = MUX_s_1_2_2(or_155_cse, exit_COMPUTE_LOOP_lpi_1_dfm_1,
      or_dcpl_63);
  assign exit_COMPUTE_LOOP_lpi_1_dfm_3_mx0w0 = COMPUTE_LOOP_mux_4_nl & exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0;
  assign CONVOLUTION_LOOP_mux_1_nl = MUX_s_1_2_2(or_157_cse, exit_CONVOLUTION_LOOP_lpi_1_dfm_1,
      or_dcpl_62);
  assign exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0 = CONVOLUTION_LOOP_mux_1_nl & exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0w0;
  assign exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0 = exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0
      & main_stage_v_1;
  assign CONVOLUTION_LOOP_for_mux_6_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_sva_2_mx0w0,
      exit_CONVOLUTION_LOOP_for_sva_2, or_dcpl_76);
  assign exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0w0 = ((CONVOLUTION_LOOP_for_acc_tmp[5])
      | CONVOLUTION_LOOP_for_mux_6_nl) & exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_2_mx0w0;
  assign exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0 = exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0w0
      & main_stage_v_1;
  assign exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_2_mx0w0 = nand_52_cse & exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0;
  assign exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0 = nand_74_cse & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_4;
  assign exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1 = (exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0
      & main_stage_v_1) | exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1;
  assign exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1 = (exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_2_mx0w0
      & main_stage_v_1) | (~((~ exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0) & lfst_exit_CONVOLUTION_LOOP_1_lpi_1_dfm_1));
  assign lfst_exit_CONVOLUTION_LOOP_1_lpi_1_dfm_1 = ~(exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0
      | exitL_exit_COMPUTE_LOOP_sva_mx0);
  assign unequal_tmp_1 = ~((conf_info_rsci_idat_mxwt[7:0]==8'b00000001));
  assign nl_if_acc_4_cse_1 = ({(pad_sva_1[6:0]) , 1'b0}) - (conf_info_rsci_idat_mxwt[31:24]);
  assign if_acc_4_cse_1 = nl_if_acc_4_cse_1[7:0];
  assign operator_43_true_and_nl = (pad_acc_psp_sva_1[16]) & (pad_acc_psp_sva_1[0]);
  assign nl_operator_43_true_operator_43_true_acc_nl = (pad_acc_psp_sva_1[8:1]) +
      conv_u2s_1_8(operator_43_true_and_nl);
  assign operator_43_true_operator_43_true_acc_nl = nl_operator_43_true_operator_43_true_acc_nl[7:0];
  assign nl_pad_sva_1 = $signed(operator_43_true_operator_43_true_acc_nl) * $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[15:8]));
  assign pad_sva_1 = nl_pad_sva_1[7:0];
  assign nl_else_acc_2_psp_sva_1 = conv_u2s_10_11(else_acc_4_cse_1) + conv_s2s_9_11({1'b1
      , (conf_info_rsci_idat_mxwt[47:40])});
  assign else_acc_2_psp_sva_1 = nl_else_acc_2_psp_sva_1[10:0];
  assign nl_else_acc_4_cse_1 = conv_u2u_9_10({pad_sva_1 , 1'b0}) + conv_u2u_8_10(~
      (conf_info_rsci_idat_mxwt[31:24])) + 10'b0000000001;
  assign else_acc_4_cse_1 = nl_else_acc_4_cse_1[9:0];
  assign nl_else_acc_psp_sva_1 = conv_u2s_10_11(else_acc_4_cse_1) + conv_s2s_9_11({1'b1
      , (conf_info_rsci_idat_mxwt[55:48])});
  assign else_acc_psp_sva_1 = nl_else_acc_psp_sva_1[10:0];
  assign nl_pad_acc_2_nl = ({1'b1 , (~ (conf_info_rsci_idat_mxwt[55:48]))}) + conv_u2s_8_9(conf_info_rsci_idat_mxwt[31:24])
      + 9'b000000001;
  assign pad_acc_2_nl = nl_pad_acc_2_nl[8:0];
  assign nl_operator_8_false_acc_nl = conv_u2s_8_9(conf_info_rsci_idat_mxwt[55:48])
      + 9'b111111111;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[8:0];
  assign nl_pad_mul_nl = $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[7:0])) * $signed(operator_8_false_acc_nl);
  assign pad_mul_nl = nl_pad_mul_nl[16:0];
  assign nl_pad_acc_psp_sva_1 = conv_s2s_9_17(pad_acc_2_nl) + pad_mul_nl;
  assign pad_acc_psp_sva_1 = nl_pad_acc_psp_sva_1[16:0];
  assign conf_info_crt_lpi_1_dfm_7_0_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_7_0,
      (conf_info_rsci_idat_mxwt[7:0]), exitL_exit_COMPUTE_LOOP_sva);
  assign nl_operator_8_false_1_acc_imod_2_sva_1 = ({1'b1 , (operator_8_false_1_acc_imod_1_sva_1[0])})
      + conv_u2s_1_2(~ (operator_8_false_1_acc_imod_1_sva_1[1])) + conv_u2s_1_2(~
      (operator_8_false_1_acc_imod_1_sva_1[2]));
  assign operator_8_false_1_acc_imod_2_sva_1 = nl_operator_8_false_1_acc_imod_2_sva_1[1:0];
  assign nl_operator_8_false_1_acc_8_nl = conv_s2s_1_2(~ (operator_8_false_1_acc_imod_sva_1[3]))
      + conv_u2s_1_2(operator_8_false_1_acc_imod_sva_1[0]);
  assign operator_8_false_1_acc_8_nl = nl_operator_8_false_1_acc_8_nl[1:0];
  assign nl_operator_8_false_1_acc_7_nl = conv_u2u_1_2(~ (operator_8_false_1_acc_imod_sva_1[1]))
      + conv_u2u_1_2(operator_8_false_1_acc_imod_sva_1[2]);
  assign operator_8_false_1_acc_7_nl = nl_operator_8_false_1_acc_7_nl[1:0];
  assign nl_operator_8_false_1_acc_imod_1_sva_1 = conv_s2s_2_3(operator_8_false_1_acc_8_nl)
      + conv_u2s_2_3(operator_8_false_1_acc_7_nl);
  assign operator_8_false_1_acc_imod_1_sva_1 = nl_operator_8_false_1_acc_imod_1_sva_1[2:0];
  assign nl_operator_8_false_1_acc_4_nl = conv_u2u_1_2(~ (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[3]))
      + conv_u2u_1_2(CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[4]) + conv_u2u_1_2(~
      (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[5]));
  assign operator_8_false_1_acc_4_nl = nl_operator_8_false_1_acc_4_nl[1:0];
  assign nl_operator_8_false_1_acc_6_nl = conv_u2u_2_3(z_out_1) + conv_u2u_2_3(operator_8_false_1_acc_4_nl)
      + conv_u2u_1_3(~ (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[7]));
  assign operator_8_false_1_acc_6_nl = nl_operator_8_false_1_acc_6_nl[2:0];
  assign nl_operator_8_false_1_acc_imod_sva_1 = conv_u2s_3_4(operator_8_false_1_acc_6_nl)
      + conv_s2s_3_4({2'b10 , (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[0])});
  assign operator_8_false_1_acc_imod_sva_1 = nl_operator_8_false_1_acc_imod_sva_1[3:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_asn_2929_mx0w0 = CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1
      * conf_info_crt_lpi_1_dfm_7_0_mx0;
  assign CONVOLUTION_LOOP_for_for_for_for_asn_2929_mx0w0 = nl_CONVOLUTION_LOOP_for_for_for_for_asn_2929_mx0w0[7:0];
  assign CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0 = MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_x_lpi_1,
      CONVOLUTION_LOOP_for_for_for_for_asn_2929_mx0w0, exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1);
  assign nl_operator_8_false_2_acc_psp_1 = (operator_8_false_2_acc_5_sdt_1[3:1])
      + 3'b101;
  assign operator_8_false_2_acc_psp_1 = nl_operator_8_false_2_acc_psp_1[2:0];
  assign nl_operator_8_false_2_acc_5_sdt_1 = conv_u2u_3_4(z_out) + conv_u2u_2_4(CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[5:4])
      + conv_u2u_2_4(~ (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[7:6]));
  assign operator_8_false_2_acc_5_sdt_1 = nl_operator_8_false_2_acc_5_sdt_1[3:0];
  assign nl_operator_8_false_3_acc_4_nl = ({2'b10 , (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[1:0])})
      + conv_u2s_3_4(z_out);
  assign operator_8_false_3_acc_4_nl = nl_operator_8_false_3_acc_4_nl[3:0];
  assign nl_operator_8_false_3_acc_imod_sva_1 = conv_s2s_4_5(operator_8_false_3_acc_4_nl)
      + conv_u2s_4_5({z_out_1 , 1'b0 , (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[5])});
  assign operator_8_false_3_acc_imod_sva_1 = nl_operator_8_false_3_acc_imod_sva_1[4:0];
  assign nl_COMPUTE_LOOP_acc_tmp = conv_u2u_4_5(COMPUTE_LOOP_b_4_0_lpi_1_dfm_1_3_0)
      + 5'b00001;
  assign COMPUTE_LOOP_acc_tmp = nl_COMPUTE_LOOP_acc_tmp[4:0];
  assign nl_operator_8_false_8_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_231_224_mx0)
      + 9'b111111111;
  assign operator_8_false_8_acc_tmp = nl_operator_8_false_8_acc_tmp[8:0];
  assign conf_info_crt_lpi_1_dfm_231_224_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_231_224,
      (conf_info_rsci_idat_mxwt[63:56]), exitL_exit_COMPUTE_LOOP_sva);
  assign nl_CONVOLUTION_LOOP_acc_tmp = conv_u2u_5_6(CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_1_4_0)
      + 6'b000001;
  assign CONVOLUTION_LOOP_acc_tmp = nl_CONVOLUTION_LOOP_acc_tmp[5:0];
  assign exit_CONVOLUTION_LOOP_sva_3 = ~((~((CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_1_4_0
      == (operator_8_false_7_acc_tmp[4:0])) & (operator_8_false_7_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_7_acc_tmp[8]));
  assign nl_operator_8_false_7_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_71_64_mx0)
      + 9'b111111111;
  assign operator_8_false_7_acc_tmp = nl_operator_8_false_7_acc_tmp[8:0];
  assign conf_info_crt_lpi_1_dfm_71_64_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_71_64,
      (conf_info_rsci_idat_mxwt[23:16]), exitL_exit_COMPUTE_LOOP_sva);
  assign nl_CONVOLUTION_LOOP_for_acc_tmp = conv_u2u_5_6(CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0)
      + 6'b000001;
  assign CONVOLUTION_LOOP_for_acc_tmp = nl_CONVOLUTION_LOOP_for_acc_tmp[5:0];
  assign CONVOLUTION_LOOP_for_if_equal_tmp = CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0
      == (operator_8_false_3_acc_tmp[4:0]);
  assign exit_CONVOLUTION_LOOP_for_sva_2_mx0w0 = ~((~(CONVOLUTION_LOOP_for_if_equal_tmp
      & (operator_8_false_3_acc_tmp[7:5]==3'b000))) | (operator_8_false_3_acc_tmp[8]));
  assign CONVOLUTION_LOOP_for_for_if_CONVOLUTION_LOOP_for_for_if_nand_tmp = ~((CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1
      == (operator_8_false_5_acc_tmp[4:0])) & (operator_8_false_5_acc_tmp[7:5]==3'b000));
  assign nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2 = CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1
      + 5'b00001;
  assign CONVOLUTION_LOOP_for_for_i_4_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2[4:0];
  assign nl_operator_8_false_5_acc_tmp = conv_u2s_8_9(n_w_out_lpi_1_dfm_2) + 9'b111111111;
  assign operator_8_false_5_acc_tmp = nl_operator_8_false_5_acc_tmp[8:0];
  assign COMPUTE_LOOP_or_2_cse = ((~ unequal_tmp_1) & exitL_exit_COMPUTE_LOOP_sva)
      | (unequal_tmp_1 & exitL_exit_COMPUTE_LOOP_sva);
  assign if_mux_4_nl = MUX_v_8_2_2(if_acc_4_cse_1, (else_acc_psp_sva_1[8:1]), or_314_cse);
  assign operator_42_true_and_1_nl = (else_acc_psp_sva_1[10]) & (else_acc_psp_sva_1[0]);
  assign if_mux_5_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[55:48]), ({7'b0000000
      , operator_42_true_and_1_nl}), or_314_cse);
  assign nl_acc_3_nl = ({if_mux_4_nl , 1'b1}) + ({if_mux_5_nl , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[8:0];
  assign n_w_out_lpi_1_dfm_2 = MUX_v_8_2_2(n_w_out_lpi_1_dfm_1, (readslicef_9_8_1(acc_3_nl)),
      COMPUTE_LOOP_or_2_cse);
  assign CONVOLUTION_LOOP_for_for_for_acc_0_sva_2 = ~((~((CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1[0])
      | CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl = ~(MUX_v_55_2_2((CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1[55:1]),
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2 = ~(MUX_v_55_2_2(CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl,
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_acc_56_sva_2 = ~((~((CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1[56])
      | CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_67_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_66_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_65_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_64_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_63_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_62_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_61_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_60_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_59_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_58_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_57_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_56_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_56_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_57_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_58_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_59_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_60_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_61_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_62_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_63_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_64_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_65_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_66_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_7_67_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_67_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_66_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_65_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_64_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_63_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_62_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_61_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_60_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_59_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_58_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_57_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_56_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_55_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_54_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_53_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_52_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_51_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_50_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_49_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_48_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_47_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_46_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_45_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_44_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_43_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_42_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_41_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_40_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_39_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_38_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_37_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_36_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_35_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_32_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_34_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_33_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:3]==2'b01);
  assign nl_CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1 = conv_u2u_2_5(CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[4:3])
      + CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1;
  assign CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1 = nl_CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:0];
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_67_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_66_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_65_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_64_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_63_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_63_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_62_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_62_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_61_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_61_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_60_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_60_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_59_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_59_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_58_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_58_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_57_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_57_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_56_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_56_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_55_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_55_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_54_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_54_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_53_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_53_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_52_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_52_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_51_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_51_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_50_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_50_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_49_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_49_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_48_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_48_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_47_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_47_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_46_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_46_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_45_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_45_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_44_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_44_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_43_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_43_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_42_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_42_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_41_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_41_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_40_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_40_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_6_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_40_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_41_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_42_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_43_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_44_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_45_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_46_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_47_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_48_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_49_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_50_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_51_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_52_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_53_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_54_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_55_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_56_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_57_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_58_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_59_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_60_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_61_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_62_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_63_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_5_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1 = CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1
      + conv_u2u_4_5(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[4:1]);
  assign CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1 = nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[4:0];
  assign CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1 = ~((~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[0])
      | CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_nor_1_nl = ~(MUX_v_55_2_2((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[55:1]),
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1 = ~(MUX_v_55_2_2(CONVOLUTION_LOOP_for_for_for_else_nor_1_nl,
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1 = ~((~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[56])
      | CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_67_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_67_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_66_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_66_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_65_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_65_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_64_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_64_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_63_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_63_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_62_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_62_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_61_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_61_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_60_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_60_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_59_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_59_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_58_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_58_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_57_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_57_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_if_and_stg_7_56_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_56_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_55_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_54_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_53_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_52_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_51_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_50_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_49_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_48_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_47_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_46_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_45_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_44_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_43_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_42_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_41_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_40_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_39_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_38_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_37_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_36_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_35_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_32_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_34_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_6_33_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_63_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_62_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_61_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_60_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_59_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_58_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_57_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_56_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_55_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_54_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_53_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_52_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_51_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_50_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_49_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_48_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_47_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_46_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_45_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_44_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_43_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_42_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_41_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_40_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1 = CONVOLUTION_LOOP_for_for_for_if_and_stg_5_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])
      | (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1 = (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])
      & (~ (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1 = (~ (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0]))
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1 = (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])
      & (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_nl = MUX_s_1_324_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1, {CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1
      , (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0]) , (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])});
  assign CONVOLUTION_LOOP_for_for_for_else_mux_972_nl = MUX_v_55_324_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1, {CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1
      , (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0]) , (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])});
  assign CONVOLUTION_LOOP_for_for_for_else_mux_973_nl = MUX_s_1_324_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1, COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1,
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1, {CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1
      , (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0]) , (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])});
  assign nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1 = conv_s2s_57_58({CONVOLUTION_LOOP_for_for_for_else_mux_nl
      , CONVOLUTION_LOOP_for_for_for_else_mux_972_nl , CONVOLUTION_LOOP_for_for_for_else_mux_973_nl})
      + conv_s2s_57_58({CONVOLUTION_LOOP_for_for_for_acc_56_sva_2 , CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2
      , CONVOLUTION_LOOP_for_for_for_acc_0_sva_2});
  assign CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:0];
  assign CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:56]==2'b10);
  assign CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:56]!=2'b01));
  assign CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_55_1_1
      = MUX_v_55_324_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1_dfm_2,
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1_dfm_2, COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1_dfm_2,
      {CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1 , (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0])
      , (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])});
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1 = CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_56_1
      & (~((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_55_1_1[54:30]==25'b1111111111111111111111111)));
  assign CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1 = ~(CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_56_1
      | (~((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_55_1_1[54:30]!=25'b0000000000000000000000000))));
  assign CONVOLUTION_LOOP_for_for_for_else_mux_974_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_972_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_974_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_972_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_976_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_973_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_976_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_973_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_978_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_974_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_978_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_974_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_980_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_975_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_980_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_975_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_982_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_976_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_982_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_976_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_984_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_977_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_984_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_977_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_986_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_978_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_986_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_978_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_988_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_979_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_988_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_979_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_990_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_980_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_990_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_980_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_992_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_981_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_992_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_981_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_994_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_982_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_994_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_982_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_996_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_983_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_996_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_983_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_998_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_984_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_998_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_984_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_985_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_985_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_986_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_986_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_987_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_987_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_988_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_988_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_989_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_989_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_990_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_990_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_991_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_991_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_992_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_992_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_993_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_993_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_994_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_994_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_995_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_995_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_996_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_996_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_997_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_997_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_998_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_998_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_999_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_999_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_56_1
      = MUX_s_1_324_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1_dfm_1_mx0,
      {CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1 , (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0])
      , (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])});
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1297_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1297_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1626_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1298_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1626_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1298_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1628_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1299_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1628_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1299_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1630_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1300_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1630_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1300_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1632_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1301_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1632_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1301_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1634_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1302_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1634_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1302_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1636_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1303_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1636_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1303_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1638_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1304_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1638_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1304_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1640_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1305_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1640_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1305_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1642_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1306_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1642_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1306_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1644_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1307_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1644_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1307_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1646_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1308_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1646_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1308_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1648_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1309_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1648_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1309_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1650_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1310_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1650_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1310_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1652_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1311_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1652_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1311_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1654_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1312_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1654_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1312_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1656_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1313_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1656_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1313_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1658_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1314_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1658_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1314_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1660_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1315_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1660_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1315_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1662_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1316_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1662_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1316_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1664_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1317_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1664_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1317_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1666_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1318_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1666_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1318_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1668_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1319_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1668_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1319_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1670_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1320_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1670_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1320_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1672_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1321_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1672_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1321_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1674_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1322_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1674_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1322_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1676_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1323_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1676_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1323_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1678_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1324_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1678_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1324_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1680_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1325_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1680_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1325_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1682_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1326_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1682_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1326_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1684_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1327_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1684_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1327_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1686_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1328_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1686_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1328_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1688_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1329_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1688_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1329_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1690_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1330_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1690_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1330_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1692_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1331_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1692_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1331_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1694_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1332_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1694_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1332_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1696_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1333_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1696_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1333_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1698_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1334_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1698_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1334_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1700_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1335_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1700_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1335_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1702_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1336_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1702_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1336_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1704_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1337_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1704_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1337_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1706_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1338_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1706_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1338_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1708_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1339_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1708_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1339_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1710_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1340_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1710_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1340_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1712_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1341_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1712_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1341_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1714_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1342_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1714_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1342_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1716_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1343_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1716_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1343_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1718_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1344_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1718_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1344_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1720_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1345_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1720_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1345_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1722_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1346_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1722_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1346_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1724_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1347_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1724_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1347_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1726_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1348_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1726_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1348_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1728_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1349_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1728_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1349_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1730_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1350_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1730_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1350_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1732_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1351_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1732_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1351_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1734_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1352_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1734_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1352_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1736_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1353_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1736_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1353_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1738_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1354_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1738_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1354_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1740_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1355_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1740_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1355_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1742_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1356_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1742_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1356_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1744_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1357_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1744_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1357_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1746_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1358_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1746_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1358_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1748_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1359_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1748_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1359_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1750_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1360_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1750_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1360_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1752_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1361_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1752_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1361_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1754_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1362_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1754_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1362_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1756_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1363_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1756_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1363_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1758_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1364_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1758_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1364_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1760_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1365_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1760_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1365_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1762_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1366_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1762_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1366_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1764_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1367_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1764_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1367_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1766_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1368_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1766_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1368_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1768_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1369_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1768_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1369_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1770_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1370_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1770_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1370_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1772_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1371_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1772_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1371_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1774_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1372_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1774_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1372_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1776_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1373_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1776_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1373_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1778_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1374_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1778_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1374_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1780_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1375_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1780_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1375_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1782_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1376_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1782_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1376_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1784_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1377_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1784_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1377_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1786_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1378_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1786_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1378_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1788_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1379_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1788_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1379_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1790_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1380_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1790_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1380_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1792_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1381_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1792_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1381_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1794_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1382_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1794_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1382_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1796_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1383_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1796_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1383_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1798_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1384_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1798_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1384_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1800_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1385_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1800_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1385_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1802_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1386_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1802_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1386_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1804_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1387_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1804_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1387_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1806_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1388_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1806_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1388_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1808_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1389_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1808_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1389_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1810_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1390_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1810_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1390_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1812_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1391_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1812_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1391_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1814_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1392_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1814_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1392_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1816_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1393_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1816_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1393_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1818_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1394_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1818_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1394_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1820_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1395_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1820_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1395_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1822_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1396_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1822_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1396_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1824_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1397_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1824_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1397_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1826_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1398_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1826_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1398_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1828_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1399_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1828_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1399_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1830_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1400_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1830_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1400_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1832_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1401_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1832_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1401_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1834_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1402_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1834_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1402_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1836_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1403_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1836_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1403_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1838_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1404_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1838_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1404_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1840_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1405_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1840_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1405_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1842_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1406_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1842_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1406_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1844_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1407_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1844_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1407_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1846_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1408_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1846_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1408_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1848_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1409_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1848_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1409_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1850_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1410_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1850_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1410_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1852_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1411_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1852_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1411_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1854_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1412_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1854_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1412_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1856_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1413_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1856_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1413_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1858_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1414_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1858_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1414_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1860_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1415_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1860_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1415_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1862_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1416_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1862_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1416_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1864_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1417_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1864_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1417_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1866_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1418_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1866_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1418_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1868_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1419_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1868_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1419_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1870_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1420_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1870_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1420_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1872_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1421_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1872_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1421_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1874_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1422_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1874_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1422_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1876_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1423_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1876_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1423_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1878_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1424_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1878_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1424_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1880_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1425_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1880_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1425_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1882_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1426_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1882_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1426_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1884_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1427_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1884_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1427_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1886_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1428_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1886_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1428_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1888_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1429_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1888_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1429_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1890_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1430_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1890_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1430_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1892_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1431_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1892_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1431_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1894_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1432_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1894_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1432_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1896_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1433_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1896_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1433_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1898_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1434_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1898_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1434_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1900_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1435_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1900_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1435_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1902_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1436_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1902_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1436_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1904_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1437_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1904_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1437_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1906_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1438_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1906_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1438_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1908_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1439_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1908_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1439_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1910_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1440_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1910_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1440_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1912_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1441_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1912_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1441_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1914_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1442_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1914_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1442_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1916_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1443_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1916_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1443_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1918_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1444_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1918_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1444_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1920_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1445_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1920_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1445_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1922_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1446_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1922_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1446_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1924_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1447_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1924_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1447_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1926_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1448_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1926_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1448_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1928_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1449_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1928_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1449_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1930_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1450_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1930_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1450_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1932_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1451_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1932_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1451_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1934_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1452_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1934_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1452_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1936_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1453_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1936_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1453_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1938_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1454_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1938_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1454_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1940_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1455_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1940_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1455_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1942_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1456_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1942_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1456_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1944_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1457_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1944_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1457_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1946_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1458_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1946_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1458_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1948_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1459_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1948_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1459_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1950_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1460_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1950_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1460_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1952_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1461_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1952_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1461_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1954_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1462_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1954_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1462_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1956_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1463_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1956_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1463_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1958_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1464_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1958_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1464_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1960_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1465_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1960_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1465_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1962_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1466_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1962_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1466_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1964_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1467_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1964_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1467_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1966_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1468_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1966_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1468_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1968_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1469_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1968_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1469_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1970_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1470_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1970_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1470_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1972_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1471_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1972_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1471_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1974_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1472_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1974_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1472_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1976_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1473_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1976_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1473_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1978_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1474_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1978_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1474_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1980_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1475_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1980_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1475_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1982_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1476_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1982_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1476_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1984_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1477_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1984_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1477_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1986_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1478_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1986_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1478_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1988_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1479_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1988_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1479_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1990_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1480_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1990_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1480_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1992_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1481_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1992_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1481_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1994_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1482_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1994_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1482_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1996_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1483_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1996_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1483_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1998_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1484_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_1998_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1484_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2000_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1485_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2000_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1485_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2002_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1486_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2002_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1486_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2004_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1487_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2004_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1487_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2006_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1488_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2006_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1488_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2008_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1489_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2008_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1489_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2010_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1490_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2010_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1490_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2012_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1491_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2012_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1491_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2014_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1492_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2014_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1492_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2016_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1493_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2016_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1493_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2018_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1494_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2018_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1494_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2020_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1495_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2020_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1495_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2022_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1496_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2022_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1496_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2024_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1497_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2024_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1497_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2026_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1498_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2026_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1498_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2028_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1499_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2028_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1499_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2030_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1500_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2030_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1500_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2032_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1501_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2032_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1501_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2034_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1502_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2034_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1502_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2036_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1503_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2036_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1503_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2038_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1504_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2038_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1504_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2040_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1505_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2040_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1505_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2042_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1506_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2042_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1506_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2044_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1507_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2044_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1507_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2046_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1508_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2046_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1508_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2048_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1509_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2048_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1509_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2050_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1510_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2050_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1510_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2052_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1511_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2052_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1511_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2054_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1512_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2054_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1512_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2056_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1513_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2056_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1513_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2058_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1514_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2058_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1514_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2060_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1515_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2060_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1515_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2062_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1516_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2062_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1516_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2064_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1517_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2064_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1517_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2066_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1518_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2066_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1518_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2068_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1519_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2068_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1519_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2070_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1520_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2070_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1520_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2072_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1521_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2072_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1521_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2074_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1522_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2074_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1522_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2076_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1523_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2076_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1523_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2078_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1524_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2078_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1524_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2080_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1525_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2080_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1525_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2082_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1526_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2082_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1526_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2084_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1527_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2084_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1527_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2086_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1528_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2086_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1528_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2088_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1529_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2088_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1529_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2090_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1530_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2090_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1530_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2092_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1531_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2092_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1531_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2094_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1532_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2094_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1532_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2096_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1533_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2096_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1533_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2098_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1534_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2098_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1534_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2100_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1535_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2100_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1535_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2102_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1536_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2102_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1536_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2104_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1537_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2104_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1537_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2106_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1538_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2106_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1538_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2108_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1539_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2108_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1539_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2110_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1540_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2110_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1540_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2112_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1541_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2112_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1541_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2114_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1542_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2114_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1542_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2116_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1543_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2116_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1543_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2118_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1544_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2118_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1544_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2120_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1545_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2120_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1545_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2122_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1546_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2122_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1546_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2124_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1547_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2124_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1547_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2126_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1548_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2126_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1548_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2128_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1549_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2128_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1549_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2130_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1550_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2130_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1550_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2132_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1551_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2132_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1551_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2134_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1552_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2134_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1552_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2136_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1553_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2136_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1553_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2138_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1554_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2138_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1554_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2140_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1555_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2140_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1555_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2142_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1556_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2142_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1556_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2144_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1557_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2144_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1557_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2146_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1558_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2146_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1558_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2148_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1559_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2148_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1559_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2150_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1560_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2150_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1560_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2152_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1561_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2152_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1561_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2154_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1562_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2154_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1562_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2156_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1563_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2156_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1563_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2158_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1564_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2158_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1564_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2160_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1565_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2160_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1565_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2162_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1566_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2162_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1566_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2164_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1567_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2164_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1567_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2166_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1568_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2166_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1568_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2168_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1569_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2168_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1569_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2170_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1570_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2170_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1570_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2172_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1571_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2172_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1571_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2174_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1572_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2174_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1572_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2176_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1573_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2176_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1573_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2178_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1574_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2178_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1574_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2180_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1575_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2180_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1575_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2182_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1576_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2182_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1576_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2184_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1577_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2184_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1577_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2186_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1578_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2186_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1578_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2188_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1579_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2188_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1579_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2190_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1580_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2190_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1580_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2192_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1581_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2192_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1581_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2194_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1582_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2194_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1582_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2196_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1583_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2196_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1583_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2198_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1584_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2198_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1584_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2200_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1585_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2200_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1585_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2202_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1586_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2202_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1586_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2204_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1587_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2204_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1587_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2206_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1588_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2206_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1588_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2208_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1589_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2208_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1589_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2210_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1590_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2210_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1590_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2212_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1591_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2212_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1591_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2214_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1592_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2214_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1592_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2216_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1593_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2216_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1593_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2218_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1594_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2218_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1594_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2220_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1595_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2220_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1595_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2222_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1596_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2222_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1596_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2224_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1597_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2224_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1597_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2226_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1598_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2226_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1598_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2228_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1599_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2228_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1599_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2230_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1600_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2230_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1600_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2232_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1601_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2232_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1601_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2234_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1602_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2234_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1602_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2236_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1603_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2236_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1603_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2238_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1604_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2238_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1604_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2240_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1605_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2240_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1605_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2242_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1606_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2242_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1606_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2244_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1607_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2244_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1607_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2246_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1608_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2246_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1608_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2248_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1609_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2248_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1609_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2250_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1610_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2250_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1610_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2252_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1611_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2252_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1611_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2254_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1612_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2254_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1612_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2256_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1613_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2256_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1613_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2258_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1614_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2258_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1614_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2260_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1615_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2260_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1615_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2262_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1616_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2262_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1616_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2264_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1617_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2264_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1617_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2266_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1618_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2266_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1618_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_2268_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1619_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_56_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_2268_nl,
      CONVOLUTION_LOOP_for_for_for_if_mux_1619_nl, and_dcpl_61);
  assign CONVOLUTION_LOOP_for_for_for_or_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_2_nl = CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_3_nl = CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_nl , CONVOLUTION_LOOP_for_for_for_and_2_nl
      , CONVOLUTION_LOOP_for_for_for_and_3_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_1_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_6_nl = CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_7_nl = CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_1_nl , CONVOLUTION_LOOP_for_for_for_and_6_nl
      , CONVOLUTION_LOOP_for_for_for_and_7_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_2_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_10_nl = CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_11_nl = CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_2_nl , CONVOLUTION_LOOP_for_for_for_and_10_nl
      , CONVOLUTION_LOOP_for_for_for_and_11_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_3_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_14_nl = CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_15_nl = CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_3_nl , CONVOLUTION_LOOP_for_for_for_and_14_nl
      , CONVOLUTION_LOOP_for_for_for_and_15_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_4_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_18_nl = CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_19_nl = CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_4_nl , CONVOLUTION_LOOP_for_for_for_and_18_nl
      , CONVOLUTION_LOOP_for_for_for_and_19_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_5_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_22_nl = CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_23_nl = CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_5_nl , CONVOLUTION_LOOP_for_for_for_and_22_nl
      , CONVOLUTION_LOOP_for_for_for_and_23_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_6_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_26_nl = CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_27_nl = CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_6_nl , CONVOLUTION_LOOP_for_for_for_and_26_nl
      , CONVOLUTION_LOOP_for_for_for_and_27_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_7_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_30_nl = CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_31_nl = CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_7_nl , CONVOLUTION_LOOP_for_for_for_and_30_nl
      , CONVOLUTION_LOOP_for_for_for_and_31_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_8_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_34_nl = CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_35_nl = CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_8_nl , CONVOLUTION_LOOP_for_for_for_and_34_nl
      , CONVOLUTION_LOOP_for_for_for_and_35_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_9_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_38_nl = CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_39_nl = CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_9_nl , CONVOLUTION_LOOP_for_for_for_and_38_nl
      , CONVOLUTION_LOOP_for_for_for_and_39_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_10_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_42_nl = CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_43_nl = CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_10_nl , CONVOLUTION_LOOP_for_for_for_and_42_nl
      , CONVOLUTION_LOOP_for_for_for_and_43_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_11_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_46_nl = CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_47_nl = CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_11_nl , CONVOLUTION_LOOP_for_for_for_and_46_nl
      , CONVOLUTION_LOOP_for_for_for_and_47_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_12_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_50_nl = CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_51_nl = CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_12_nl , CONVOLUTION_LOOP_for_for_for_and_50_nl
      , CONVOLUTION_LOOP_for_for_for_and_51_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_13_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_54_nl = CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_55_nl = CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_13_nl , CONVOLUTION_LOOP_for_for_for_and_54_nl
      , CONVOLUTION_LOOP_for_for_for_and_55_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_14_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_58_nl = CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_59_nl = CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_14_nl , CONVOLUTION_LOOP_for_for_for_and_58_nl
      , CONVOLUTION_LOOP_for_for_for_and_59_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_15_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_62_nl = CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_63_nl = CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_15_nl , CONVOLUTION_LOOP_for_for_for_and_62_nl
      , CONVOLUTION_LOOP_for_for_for_and_63_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_16_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_66_nl = CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_67_nl = CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_16_nl , CONVOLUTION_LOOP_for_for_for_and_66_nl
      , CONVOLUTION_LOOP_for_for_for_and_67_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_17_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_70_nl = CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_71_nl = CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_17_nl , CONVOLUTION_LOOP_for_for_for_and_70_nl
      , CONVOLUTION_LOOP_for_for_for_and_71_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_18_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_74_nl = CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_75_nl = CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_18_nl , CONVOLUTION_LOOP_for_for_for_and_74_nl
      , CONVOLUTION_LOOP_for_for_for_and_75_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_19_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_78_nl = CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_79_nl = CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_19_nl , CONVOLUTION_LOOP_for_for_for_and_78_nl
      , CONVOLUTION_LOOP_for_for_for_and_79_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_20_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_82_nl = CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_83_nl = CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_20_nl , CONVOLUTION_LOOP_for_for_for_and_82_nl
      , CONVOLUTION_LOOP_for_for_for_and_83_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_21_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_86_nl = CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_87_nl = CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_21_nl , CONVOLUTION_LOOP_for_for_for_and_86_nl
      , CONVOLUTION_LOOP_for_for_for_and_87_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_22_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_90_nl = CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_91_nl = CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_22_nl , CONVOLUTION_LOOP_for_for_for_and_90_nl
      , CONVOLUTION_LOOP_for_for_for_and_91_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_23_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_94_nl = CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_95_nl = CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_23_nl , CONVOLUTION_LOOP_for_for_for_and_94_nl
      , CONVOLUTION_LOOP_for_for_for_and_95_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_24_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_98_nl = CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_99_nl = CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_24_nl , CONVOLUTION_LOOP_for_for_for_and_98_nl
      , CONVOLUTION_LOOP_for_for_for_and_99_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_25_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_102_nl = CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_103_nl = CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_25_nl , CONVOLUTION_LOOP_for_for_for_and_102_nl
      , CONVOLUTION_LOOP_for_for_for_and_103_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_26_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_106_nl = CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_107_nl = CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_26_nl , CONVOLUTION_LOOP_for_for_for_and_106_nl
      , CONVOLUTION_LOOP_for_for_for_and_107_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_27_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_110_nl = CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_111_nl = CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_27_nl , CONVOLUTION_LOOP_for_for_for_and_110_nl
      , CONVOLUTION_LOOP_for_for_for_and_111_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_28_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_114_nl = CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_115_nl = CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_28_nl , CONVOLUTION_LOOP_for_for_for_and_114_nl
      , CONVOLUTION_LOOP_for_for_for_and_115_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_29_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_118_nl = CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_119_nl = CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_29_nl , CONVOLUTION_LOOP_for_for_for_and_118_nl
      , CONVOLUTION_LOOP_for_for_for_and_119_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_30_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_122_nl = CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_123_nl = CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_30_nl , CONVOLUTION_LOOP_for_for_for_and_122_nl
      , CONVOLUTION_LOOP_for_for_for_and_123_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_31_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_126_nl = CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_127_nl = CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_31_nl , CONVOLUTION_LOOP_for_for_for_and_126_nl
      , CONVOLUTION_LOOP_for_for_for_and_127_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_32_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_130_nl = CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_131_nl = CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_32_nl , CONVOLUTION_LOOP_for_for_for_and_130_nl
      , CONVOLUTION_LOOP_for_for_for_and_131_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_33_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_134_nl = CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_135_nl = CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_33_nl , CONVOLUTION_LOOP_for_for_for_and_134_nl
      , CONVOLUTION_LOOP_for_for_for_and_135_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_34_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_138_nl = CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_139_nl = CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_34_nl , CONVOLUTION_LOOP_for_for_for_and_138_nl
      , CONVOLUTION_LOOP_for_for_for_and_139_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_35_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_142_nl = CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_143_nl = CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_35_nl , CONVOLUTION_LOOP_for_for_for_and_142_nl
      , CONVOLUTION_LOOP_for_for_for_and_143_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_36_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_146_nl = CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_147_nl = CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_36_nl , CONVOLUTION_LOOP_for_for_for_and_146_nl
      , CONVOLUTION_LOOP_for_for_for_and_147_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_37_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_150_nl = CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_151_nl = CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_37_nl , CONVOLUTION_LOOP_for_for_for_and_150_nl
      , CONVOLUTION_LOOP_for_for_for_and_151_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_38_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_154_nl = CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_155_nl = CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_38_nl , CONVOLUTION_LOOP_for_for_for_and_154_nl
      , CONVOLUTION_LOOP_for_for_for_and_155_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_39_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_158_nl = CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_159_nl = CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_39_nl , CONVOLUTION_LOOP_for_for_for_and_158_nl
      , CONVOLUTION_LOOP_for_for_for_and_159_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_40_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_162_nl = CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_163_nl = CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_40_nl , CONVOLUTION_LOOP_for_for_for_and_162_nl
      , CONVOLUTION_LOOP_for_for_for_and_163_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_41_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_166_nl = CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_167_nl = CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_41_nl , CONVOLUTION_LOOP_for_for_for_and_166_nl
      , CONVOLUTION_LOOP_for_for_for_and_167_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_42_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_170_nl = CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_171_nl = CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_42_nl , CONVOLUTION_LOOP_for_for_for_and_170_nl
      , CONVOLUTION_LOOP_for_for_for_and_171_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_43_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_174_nl = CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_175_nl = CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_43_nl , CONVOLUTION_LOOP_for_for_for_and_174_nl
      , CONVOLUTION_LOOP_for_for_for_and_175_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_44_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_178_nl = CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_179_nl = CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_44_nl , CONVOLUTION_LOOP_for_for_for_and_178_nl
      , CONVOLUTION_LOOP_for_for_for_and_179_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_45_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_182_nl = CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_183_nl = CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_45_nl , CONVOLUTION_LOOP_for_for_for_and_182_nl
      , CONVOLUTION_LOOP_for_for_for_and_183_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_46_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_186_nl = CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_187_nl = CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_46_nl , CONVOLUTION_LOOP_for_for_for_and_186_nl
      , CONVOLUTION_LOOP_for_for_for_and_187_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_47_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_190_nl = CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_191_nl = CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_47_nl , CONVOLUTION_LOOP_for_for_for_and_190_nl
      , CONVOLUTION_LOOP_for_for_for_and_191_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_48_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_194_nl = CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_195_nl = CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_48_nl , CONVOLUTION_LOOP_for_for_for_and_194_nl
      , CONVOLUTION_LOOP_for_for_for_and_195_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_49_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_198_nl = CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_199_nl = CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_49_nl , CONVOLUTION_LOOP_for_for_for_and_198_nl
      , CONVOLUTION_LOOP_for_for_for_and_199_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_50_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_202_nl = CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_203_nl = CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_50_nl , CONVOLUTION_LOOP_for_for_for_and_202_nl
      , CONVOLUTION_LOOP_for_for_for_and_203_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_51_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_206_nl = CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_207_nl = CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_51_nl , CONVOLUTION_LOOP_for_for_for_and_206_nl
      , CONVOLUTION_LOOP_for_for_for_and_207_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_52_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_210_nl = CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_211_nl = CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_52_nl , CONVOLUTION_LOOP_for_for_for_and_210_nl
      , CONVOLUTION_LOOP_for_for_for_and_211_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_53_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_214_nl = CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_215_nl = CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_53_nl , CONVOLUTION_LOOP_for_for_for_and_214_nl
      , CONVOLUTION_LOOP_for_for_for_and_215_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_54_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_218_nl = CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_219_nl = CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_54_nl , CONVOLUTION_LOOP_for_for_for_and_218_nl
      , CONVOLUTION_LOOP_for_for_for_and_219_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_55_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_222_nl = CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_223_nl = CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_55_nl , CONVOLUTION_LOOP_for_for_for_and_222_nl
      , CONVOLUTION_LOOP_for_for_for_and_223_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_56_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_226_nl = CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_227_nl = CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_56_nl , CONVOLUTION_LOOP_for_for_for_and_226_nl
      , CONVOLUTION_LOOP_for_for_for_and_227_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_57_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_230_nl = CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_231_nl = CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_57_nl , CONVOLUTION_LOOP_for_for_for_and_230_nl
      , CONVOLUTION_LOOP_for_for_for_and_231_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_58_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_234_nl = CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_235_nl = CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_58_nl , CONVOLUTION_LOOP_for_for_for_and_234_nl
      , CONVOLUTION_LOOP_for_for_for_and_235_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_59_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_238_nl = CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_239_nl = CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_59_nl , CONVOLUTION_LOOP_for_for_for_and_238_nl
      , CONVOLUTION_LOOP_for_for_for_and_239_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_60_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_242_nl = CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_243_nl = CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_60_nl , CONVOLUTION_LOOP_for_for_for_and_242_nl
      , CONVOLUTION_LOOP_for_for_for_and_243_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_61_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_246_nl = CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_247_nl = CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_61_nl , CONVOLUTION_LOOP_for_for_for_and_246_nl
      , CONVOLUTION_LOOP_for_for_for_and_247_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_62_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_250_nl = CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_251_nl = CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_62_nl , CONVOLUTION_LOOP_for_for_for_and_250_nl
      , CONVOLUTION_LOOP_for_for_for_and_251_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_63_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_254_nl = CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_255_nl = CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_63_nl , CONVOLUTION_LOOP_for_for_for_and_254_nl
      , CONVOLUTION_LOOP_for_for_for_and_255_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_64_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_258_nl = CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_259_nl = CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_64_nl , CONVOLUTION_LOOP_for_for_for_and_258_nl
      , CONVOLUTION_LOOP_for_for_for_and_259_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_65_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_262_nl = CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_263_nl = CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_65_nl , CONVOLUTION_LOOP_for_for_for_and_262_nl
      , CONVOLUTION_LOOP_for_for_for_and_263_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_66_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_266_nl = CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_267_nl = CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_66_nl , CONVOLUTION_LOOP_for_for_for_and_266_nl
      , CONVOLUTION_LOOP_for_for_for_and_267_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_67_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_270_nl = CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_271_nl = CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_67_nl , CONVOLUTION_LOOP_for_for_for_and_270_nl
      , CONVOLUTION_LOOP_for_for_for_and_271_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_68_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_274_nl = CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_275_nl = CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_68_nl , CONVOLUTION_LOOP_for_for_for_and_274_nl
      , CONVOLUTION_LOOP_for_for_for_and_275_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_69_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_278_nl = CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_279_nl = CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_69_nl , CONVOLUTION_LOOP_for_for_for_and_278_nl
      , CONVOLUTION_LOOP_for_for_for_and_279_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_70_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_282_nl = CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_283_nl = CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_70_nl , CONVOLUTION_LOOP_for_for_for_and_282_nl
      , CONVOLUTION_LOOP_for_for_for_and_283_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_71_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_286_nl = CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_287_nl = CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_71_nl , CONVOLUTION_LOOP_for_for_for_and_286_nl
      , CONVOLUTION_LOOP_for_for_for_and_287_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_72_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_290_nl = CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_291_nl = CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_72_nl , CONVOLUTION_LOOP_for_for_for_and_290_nl
      , CONVOLUTION_LOOP_for_for_for_and_291_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_73_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_294_nl = CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_295_nl = CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_73_nl , CONVOLUTION_LOOP_for_for_for_and_294_nl
      , CONVOLUTION_LOOP_for_for_for_and_295_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_74_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_298_nl = CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_299_nl = CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_74_nl , CONVOLUTION_LOOP_for_for_for_and_298_nl
      , CONVOLUTION_LOOP_for_for_for_and_299_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_75_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_302_nl = CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_303_nl = CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_75_nl , CONVOLUTION_LOOP_for_for_for_and_302_nl
      , CONVOLUTION_LOOP_for_for_for_and_303_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_76_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_306_nl = CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_307_nl = CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_76_nl , CONVOLUTION_LOOP_for_for_for_and_306_nl
      , CONVOLUTION_LOOP_for_for_for_and_307_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_77_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_310_nl = CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_311_nl = CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_77_nl , CONVOLUTION_LOOP_for_for_for_and_310_nl
      , CONVOLUTION_LOOP_for_for_for_and_311_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_78_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_314_nl = CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_315_nl = CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_78_nl , CONVOLUTION_LOOP_for_for_for_and_314_nl
      , CONVOLUTION_LOOP_for_for_for_and_315_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_79_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_318_nl = CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_319_nl = CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_79_nl , CONVOLUTION_LOOP_for_for_for_and_318_nl
      , CONVOLUTION_LOOP_for_for_for_and_319_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_80_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_322_nl = CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_323_nl = CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_80_nl , CONVOLUTION_LOOP_for_for_for_and_322_nl
      , CONVOLUTION_LOOP_for_for_for_and_323_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_81_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_326_nl = CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_327_nl = CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_81_nl , CONVOLUTION_LOOP_for_for_for_and_326_nl
      , CONVOLUTION_LOOP_for_for_for_and_327_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_82_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_330_nl = CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_331_nl = CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_82_nl , CONVOLUTION_LOOP_for_for_for_and_330_nl
      , CONVOLUTION_LOOP_for_for_for_and_331_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_83_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_334_nl = CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_335_nl = CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_83_nl , CONVOLUTION_LOOP_for_for_for_and_334_nl
      , CONVOLUTION_LOOP_for_for_for_and_335_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_84_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_338_nl = CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_339_nl = CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_84_nl , CONVOLUTION_LOOP_for_for_for_and_338_nl
      , CONVOLUTION_LOOP_for_for_for_and_339_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_85_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_342_nl = CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_343_nl = CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_85_nl , CONVOLUTION_LOOP_for_for_for_and_342_nl
      , CONVOLUTION_LOOP_for_for_for_and_343_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_86_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_346_nl = CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_347_nl = CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_86_nl , CONVOLUTION_LOOP_for_for_for_and_346_nl
      , CONVOLUTION_LOOP_for_for_for_and_347_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_87_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_350_nl = CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_351_nl = CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_87_nl , CONVOLUTION_LOOP_for_for_for_and_350_nl
      , CONVOLUTION_LOOP_for_for_for_and_351_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_88_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_354_nl = CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_355_nl = CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_88_nl , CONVOLUTION_LOOP_for_for_for_and_354_nl
      , CONVOLUTION_LOOP_for_for_for_and_355_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_89_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_358_nl = CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_359_nl = CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_89_nl , CONVOLUTION_LOOP_for_for_for_and_358_nl
      , CONVOLUTION_LOOP_for_for_for_and_359_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_90_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_362_nl = CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_363_nl = CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_90_nl , CONVOLUTION_LOOP_for_for_for_and_362_nl
      , CONVOLUTION_LOOP_for_for_for_and_363_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_91_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_366_nl = CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_367_nl = CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_91_nl , CONVOLUTION_LOOP_for_for_for_and_366_nl
      , CONVOLUTION_LOOP_for_for_for_and_367_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_92_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_370_nl = CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_371_nl = CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_92_nl , CONVOLUTION_LOOP_for_for_for_and_370_nl
      , CONVOLUTION_LOOP_for_for_for_and_371_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_93_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_374_nl = CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_375_nl = CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_93_nl , CONVOLUTION_LOOP_for_for_for_and_374_nl
      , CONVOLUTION_LOOP_for_for_for_and_375_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_94_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_378_nl = CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_379_nl = CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_94_nl , CONVOLUTION_LOOP_for_for_for_and_378_nl
      , CONVOLUTION_LOOP_for_for_for_and_379_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_95_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_382_nl = CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_383_nl = CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_95_nl , CONVOLUTION_LOOP_for_for_for_and_382_nl
      , CONVOLUTION_LOOP_for_for_for_and_383_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_96_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_386_nl = CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_387_nl = CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_96_nl , CONVOLUTION_LOOP_for_for_for_and_386_nl
      , CONVOLUTION_LOOP_for_for_for_and_387_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_97_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_390_nl = CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_391_nl = CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_97_nl , CONVOLUTION_LOOP_for_for_for_and_390_nl
      , CONVOLUTION_LOOP_for_for_for_and_391_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_98_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_394_nl = CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_395_nl = CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_98_nl , CONVOLUTION_LOOP_for_for_for_and_394_nl
      , CONVOLUTION_LOOP_for_for_for_and_395_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_99_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_398_nl = CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_399_nl = CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_99_nl , CONVOLUTION_LOOP_for_for_for_and_398_nl
      , CONVOLUTION_LOOP_for_for_for_and_399_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_100_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_402_nl = CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_403_nl = CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_100_nl , CONVOLUTION_LOOP_for_for_for_and_402_nl
      , CONVOLUTION_LOOP_for_for_for_and_403_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_101_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_406_nl = CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_407_nl = CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_101_nl , CONVOLUTION_LOOP_for_for_for_and_406_nl
      , CONVOLUTION_LOOP_for_for_for_and_407_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_102_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_410_nl = CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_411_nl = CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_102_nl , CONVOLUTION_LOOP_for_for_for_and_410_nl
      , CONVOLUTION_LOOP_for_for_for_and_411_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_103_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_414_nl = CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_415_nl = CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_103_nl , CONVOLUTION_LOOP_for_for_for_and_414_nl
      , CONVOLUTION_LOOP_for_for_for_and_415_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_104_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_418_nl = CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_419_nl = CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_104_nl , CONVOLUTION_LOOP_for_for_for_and_418_nl
      , CONVOLUTION_LOOP_for_for_for_and_419_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_105_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_422_nl = CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_423_nl = CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_105_nl , CONVOLUTION_LOOP_for_for_for_and_422_nl
      , CONVOLUTION_LOOP_for_for_for_and_423_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_106_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_426_nl = CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_427_nl = CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_106_nl , CONVOLUTION_LOOP_for_for_for_and_426_nl
      , CONVOLUTION_LOOP_for_for_for_and_427_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_107_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_430_nl = CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_431_nl = CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_107_nl , CONVOLUTION_LOOP_for_for_for_and_430_nl
      , CONVOLUTION_LOOP_for_for_for_and_431_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_108_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_434_nl = CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_435_nl = CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_108_nl , CONVOLUTION_LOOP_for_for_for_and_434_nl
      , CONVOLUTION_LOOP_for_for_for_and_435_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_109_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_438_nl = CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_439_nl = CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_109_nl , CONVOLUTION_LOOP_for_for_for_and_438_nl
      , CONVOLUTION_LOOP_for_for_for_and_439_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_110_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_442_nl = CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_443_nl = CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_110_nl , CONVOLUTION_LOOP_for_for_for_and_442_nl
      , CONVOLUTION_LOOP_for_for_for_and_443_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_111_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_446_nl = CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_447_nl = CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_111_nl , CONVOLUTION_LOOP_for_for_for_and_446_nl
      , CONVOLUTION_LOOP_for_for_for_and_447_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_112_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_450_nl = CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_451_nl = CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_112_nl , CONVOLUTION_LOOP_for_for_for_and_450_nl
      , CONVOLUTION_LOOP_for_for_for_and_451_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_113_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_454_nl = CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_455_nl = CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_113_nl , CONVOLUTION_LOOP_for_for_for_and_454_nl
      , CONVOLUTION_LOOP_for_for_for_and_455_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_114_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_458_nl = CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_459_nl = CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_114_nl , CONVOLUTION_LOOP_for_for_for_and_458_nl
      , CONVOLUTION_LOOP_for_for_for_and_459_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_115_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_462_nl = CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_463_nl = CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_115_nl , CONVOLUTION_LOOP_for_for_for_and_462_nl
      , CONVOLUTION_LOOP_for_for_for_and_463_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_116_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_466_nl = CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_467_nl = CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_116_nl , CONVOLUTION_LOOP_for_for_for_and_466_nl
      , CONVOLUTION_LOOP_for_for_for_and_467_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_117_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_470_nl = CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_471_nl = CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_117_nl , CONVOLUTION_LOOP_for_for_for_and_470_nl
      , CONVOLUTION_LOOP_for_for_for_and_471_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_118_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_474_nl = CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_475_nl = CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_118_nl , CONVOLUTION_LOOP_for_for_for_and_474_nl
      , CONVOLUTION_LOOP_for_for_for_and_475_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_119_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_478_nl = CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_479_nl = CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_119_nl , CONVOLUTION_LOOP_for_for_for_and_478_nl
      , CONVOLUTION_LOOP_for_for_for_and_479_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_120_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_482_nl = CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_483_nl = CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_120_nl , CONVOLUTION_LOOP_for_for_for_and_482_nl
      , CONVOLUTION_LOOP_for_for_for_and_483_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_121_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_486_nl = CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_487_nl = CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_121_nl , CONVOLUTION_LOOP_for_for_for_and_486_nl
      , CONVOLUTION_LOOP_for_for_for_and_487_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_122_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_490_nl = CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_491_nl = CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_122_nl , CONVOLUTION_LOOP_for_for_for_and_490_nl
      , CONVOLUTION_LOOP_for_for_for_and_491_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_123_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_494_nl = CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_495_nl = CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_123_nl , CONVOLUTION_LOOP_for_for_for_and_494_nl
      , CONVOLUTION_LOOP_for_for_for_and_495_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_124_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_498_nl = CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_499_nl = CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_124_nl , CONVOLUTION_LOOP_for_for_for_and_498_nl
      , CONVOLUTION_LOOP_for_for_for_and_499_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_125_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_502_nl = CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_503_nl = CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_125_nl , CONVOLUTION_LOOP_for_for_for_and_502_nl
      , CONVOLUTION_LOOP_for_for_for_and_503_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_126_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_506_nl = CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_507_nl = CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_126_nl , CONVOLUTION_LOOP_for_for_for_and_506_nl
      , CONVOLUTION_LOOP_for_for_for_and_507_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_127_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_510_nl = CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_511_nl = CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_127_nl , CONVOLUTION_LOOP_for_for_for_and_510_nl
      , CONVOLUTION_LOOP_for_for_for_and_511_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_128_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_514_nl = CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_515_nl = CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_128_nl , CONVOLUTION_LOOP_for_for_for_and_514_nl
      , CONVOLUTION_LOOP_for_for_for_and_515_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_129_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_518_nl = CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_519_nl = CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_129_nl , CONVOLUTION_LOOP_for_for_for_and_518_nl
      , CONVOLUTION_LOOP_for_for_for_and_519_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_130_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_522_nl = CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_523_nl = CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_130_nl , CONVOLUTION_LOOP_for_for_for_and_522_nl
      , CONVOLUTION_LOOP_for_for_for_and_523_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_131_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_526_nl = CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_527_nl = CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_131_nl , CONVOLUTION_LOOP_for_for_for_and_526_nl
      , CONVOLUTION_LOOP_for_for_for_and_527_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_132_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_530_nl = CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_531_nl = CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_132_nl , CONVOLUTION_LOOP_for_for_for_and_530_nl
      , CONVOLUTION_LOOP_for_for_for_and_531_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_133_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_534_nl = CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_535_nl = CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_133_nl , CONVOLUTION_LOOP_for_for_for_and_534_nl
      , CONVOLUTION_LOOP_for_for_for_and_535_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_134_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_538_nl = CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_539_nl = CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_134_nl , CONVOLUTION_LOOP_for_for_for_and_538_nl
      , CONVOLUTION_LOOP_for_for_for_and_539_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_135_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_542_nl = CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_543_nl = CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_135_nl , CONVOLUTION_LOOP_for_for_for_and_542_nl
      , CONVOLUTION_LOOP_for_for_for_and_543_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_136_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_546_nl = CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_547_nl = CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_136_nl , CONVOLUTION_LOOP_for_for_for_and_546_nl
      , CONVOLUTION_LOOP_for_for_for_and_547_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_137_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_550_nl = CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_551_nl = CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_137_nl , CONVOLUTION_LOOP_for_for_for_and_550_nl
      , CONVOLUTION_LOOP_for_for_for_and_551_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_138_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_554_nl = CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_555_nl = CONVOLUTION_LOOP_for_for_for_if_and_554_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_138_nl , CONVOLUTION_LOOP_for_for_for_and_554_nl
      , CONVOLUTION_LOOP_for_for_for_and_555_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_139_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_558_nl = CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_559_nl = CONVOLUTION_LOOP_for_for_for_if_and_552_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_139_nl , CONVOLUTION_LOOP_for_for_for_and_558_nl
      , CONVOLUTION_LOOP_for_for_for_and_559_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_140_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_562_nl = CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_563_nl = CONVOLUTION_LOOP_for_for_for_if_and_550_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_140_nl , CONVOLUTION_LOOP_for_for_for_and_562_nl
      , CONVOLUTION_LOOP_for_for_for_and_563_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_141_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_566_nl = CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_567_nl = CONVOLUTION_LOOP_for_for_for_if_and_548_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_141_nl , CONVOLUTION_LOOP_for_for_for_and_566_nl
      , CONVOLUTION_LOOP_for_for_for_and_567_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_142_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_570_nl = CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_571_nl = CONVOLUTION_LOOP_for_for_for_if_and_546_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_142_nl , CONVOLUTION_LOOP_for_for_for_and_570_nl
      , CONVOLUTION_LOOP_for_for_for_and_571_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_143_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_574_nl = CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_575_nl = CONVOLUTION_LOOP_for_for_for_if_and_544_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_143_nl , CONVOLUTION_LOOP_for_for_for_and_574_nl
      , CONVOLUTION_LOOP_for_for_for_and_575_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_144_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_578_nl = CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_579_nl = CONVOLUTION_LOOP_for_for_for_if_and_542_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_144_nl , CONVOLUTION_LOOP_for_for_for_and_578_nl
      , CONVOLUTION_LOOP_for_for_for_and_579_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_145_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_582_nl = CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_583_nl = CONVOLUTION_LOOP_for_for_for_if_and_540_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_145_nl , CONVOLUTION_LOOP_for_for_for_and_582_nl
      , CONVOLUTION_LOOP_for_for_for_and_583_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_146_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_586_nl = CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_587_nl = CONVOLUTION_LOOP_for_for_for_if_and_538_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_146_nl , CONVOLUTION_LOOP_for_for_for_and_586_nl
      , CONVOLUTION_LOOP_for_for_for_and_587_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_147_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_590_nl = CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_591_nl = CONVOLUTION_LOOP_for_for_for_if_and_536_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_147_nl , CONVOLUTION_LOOP_for_for_for_and_590_nl
      , CONVOLUTION_LOOP_for_for_for_and_591_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_148_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_594_nl = CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_595_nl = CONVOLUTION_LOOP_for_for_for_if_and_534_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_148_nl , CONVOLUTION_LOOP_for_for_for_and_594_nl
      , CONVOLUTION_LOOP_for_for_for_and_595_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_149_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_598_nl = CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_599_nl = CONVOLUTION_LOOP_for_for_for_if_and_532_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_149_nl , CONVOLUTION_LOOP_for_for_for_and_598_nl
      , CONVOLUTION_LOOP_for_for_for_and_599_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_150_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_602_nl = CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_603_nl = CONVOLUTION_LOOP_for_for_for_if_and_530_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_150_nl , CONVOLUTION_LOOP_for_for_for_and_602_nl
      , CONVOLUTION_LOOP_for_for_for_and_603_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_151_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_606_nl = CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_607_nl = CONVOLUTION_LOOP_for_for_for_if_and_528_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_151_nl , CONVOLUTION_LOOP_for_for_for_and_606_nl
      , CONVOLUTION_LOOP_for_for_for_and_607_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_152_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_610_nl = CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_611_nl = CONVOLUTION_LOOP_for_for_for_if_and_526_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_152_nl , CONVOLUTION_LOOP_for_for_for_and_610_nl
      , CONVOLUTION_LOOP_for_for_for_and_611_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_153_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_614_nl = CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_615_nl = CONVOLUTION_LOOP_for_for_for_if_and_524_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_153_nl , CONVOLUTION_LOOP_for_for_for_and_614_nl
      , CONVOLUTION_LOOP_for_for_for_and_615_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_154_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_618_nl = CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_619_nl = CONVOLUTION_LOOP_for_for_for_if_and_522_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_154_nl , CONVOLUTION_LOOP_for_for_for_and_618_nl
      , CONVOLUTION_LOOP_for_for_for_and_619_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_155_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_622_nl = CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_623_nl = CONVOLUTION_LOOP_for_for_for_if_and_520_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_155_nl , CONVOLUTION_LOOP_for_for_for_and_622_nl
      , CONVOLUTION_LOOP_for_for_for_and_623_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_156_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_626_nl = CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_627_nl = CONVOLUTION_LOOP_for_for_for_if_and_518_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_156_nl , CONVOLUTION_LOOP_for_for_for_and_626_nl
      , CONVOLUTION_LOOP_for_for_for_and_627_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_157_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_630_nl = CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_631_nl = CONVOLUTION_LOOP_for_for_for_if_and_516_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_157_nl , CONVOLUTION_LOOP_for_for_for_and_630_nl
      , CONVOLUTION_LOOP_for_for_for_and_631_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_158_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_634_nl = CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_635_nl = CONVOLUTION_LOOP_for_for_for_if_and_514_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_158_nl , CONVOLUTION_LOOP_for_for_for_and_634_nl
      , CONVOLUTION_LOOP_for_for_for_and_635_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_159_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_638_nl = CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_639_nl = CONVOLUTION_LOOP_for_for_for_if_and_512_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_159_nl , CONVOLUTION_LOOP_for_for_for_and_638_nl
      , CONVOLUTION_LOOP_for_for_for_and_639_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_160_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_642_nl = CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_643_nl = CONVOLUTION_LOOP_for_for_for_if_and_510_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_160_nl , CONVOLUTION_LOOP_for_for_for_and_642_nl
      , CONVOLUTION_LOOP_for_for_for_and_643_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_161_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_646_nl = CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_647_nl = CONVOLUTION_LOOP_for_for_for_if_and_508_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_161_nl , CONVOLUTION_LOOP_for_for_for_and_646_nl
      , CONVOLUTION_LOOP_for_for_for_and_647_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_162_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_650_nl = CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_651_nl = CONVOLUTION_LOOP_for_for_for_if_and_509_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_162_nl , CONVOLUTION_LOOP_for_for_for_and_650_nl
      , CONVOLUTION_LOOP_for_for_for_and_651_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_163_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_654_nl = CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_655_nl = CONVOLUTION_LOOP_for_for_for_if_and_511_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_163_nl , CONVOLUTION_LOOP_for_for_for_and_654_nl
      , CONVOLUTION_LOOP_for_for_for_and_655_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_164_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_658_nl = CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_659_nl = CONVOLUTION_LOOP_for_for_for_if_and_513_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_164_nl , CONVOLUTION_LOOP_for_for_for_and_658_nl
      , CONVOLUTION_LOOP_for_for_for_and_659_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_165_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_662_nl = CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_663_nl = CONVOLUTION_LOOP_for_for_for_if_and_515_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_165_nl , CONVOLUTION_LOOP_for_for_for_and_662_nl
      , CONVOLUTION_LOOP_for_for_for_and_663_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_166_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_666_nl = CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_667_nl = CONVOLUTION_LOOP_for_for_for_if_and_517_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_166_nl , CONVOLUTION_LOOP_for_for_for_and_666_nl
      , CONVOLUTION_LOOP_for_for_for_and_667_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_167_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_670_nl = CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_671_nl = CONVOLUTION_LOOP_for_for_for_if_and_519_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_167_nl , CONVOLUTION_LOOP_for_for_for_and_670_nl
      , CONVOLUTION_LOOP_for_for_for_and_671_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_168_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_674_nl = CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_675_nl = CONVOLUTION_LOOP_for_for_for_if_and_521_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_168_nl , CONVOLUTION_LOOP_for_for_for_and_674_nl
      , CONVOLUTION_LOOP_for_for_for_and_675_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_169_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_678_nl = CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_679_nl = CONVOLUTION_LOOP_for_for_for_if_and_523_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_169_nl , CONVOLUTION_LOOP_for_for_for_and_678_nl
      , CONVOLUTION_LOOP_for_for_for_and_679_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_170_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_682_nl = CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_683_nl = CONVOLUTION_LOOP_for_for_for_if_and_525_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_170_nl , CONVOLUTION_LOOP_for_for_for_and_682_nl
      , CONVOLUTION_LOOP_for_for_for_and_683_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_171_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_686_nl = CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_687_nl = CONVOLUTION_LOOP_for_for_for_if_and_527_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_171_nl , CONVOLUTION_LOOP_for_for_for_and_686_nl
      , CONVOLUTION_LOOP_for_for_for_and_687_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_172_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_690_nl = CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_691_nl = CONVOLUTION_LOOP_for_for_for_if_and_529_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_172_nl , CONVOLUTION_LOOP_for_for_for_and_690_nl
      , CONVOLUTION_LOOP_for_for_for_and_691_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_173_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_694_nl = CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_695_nl = CONVOLUTION_LOOP_for_for_for_if_and_531_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_173_nl , CONVOLUTION_LOOP_for_for_for_and_694_nl
      , CONVOLUTION_LOOP_for_for_for_and_695_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_174_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_698_nl = CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_699_nl = CONVOLUTION_LOOP_for_for_for_if_and_533_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_174_nl , CONVOLUTION_LOOP_for_for_for_and_698_nl
      , CONVOLUTION_LOOP_for_for_for_and_699_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_175_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_702_nl = CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_703_nl = CONVOLUTION_LOOP_for_for_for_if_and_535_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_175_nl , CONVOLUTION_LOOP_for_for_for_and_702_nl
      , CONVOLUTION_LOOP_for_for_for_and_703_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_176_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_706_nl = CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_707_nl = CONVOLUTION_LOOP_for_for_for_if_and_537_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_176_nl , CONVOLUTION_LOOP_for_for_for_and_706_nl
      , CONVOLUTION_LOOP_for_for_for_and_707_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_177_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_710_nl = CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_711_nl = CONVOLUTION_LOOP_for_for_for_if_and_539_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_177_nl , CONVOLUTION_LOOP_for_for_for_and_710_nl
      , CONVOLUTION_LOOP_for_for_for_and_711_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_178_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_714_nl = CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_715_nl = CONVOLUTION_LOOP_for_for_for_if_and_541_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_178_nl , CONVOLUTION_LOOP_for_for_for_and_714_nl
      , CONVOLUTION_LOOP_for_for_for_and_715_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_179_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_718_nl = CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_719_nl = CONVOLUTION_LOOP_for_for_for_if_and_543_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_179_nl , CONVOLUTION_LOOP_for_for_for_and_718_nl
      , CONVOLUTION_LOOP_for_for_for_and_719_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_180_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_722_nl = CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_723_nl = CONVOLUTION_LOOP_for_for_for_if_and_545_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_180_nl , CONVOLUTION_LOOP_for_for_for_and_722_nl
      , CONVOLUTION_LOOP_for_for_for_and_723_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_181_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_726_nl = CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_727_nl = CONVOLUTION_LOOP_for_for_for_if_and_547_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_181_nl , CONVOLUTION_LOOP_for_for_for_and_726_nl
      , CONVOLUTION_LOOP_for_for_for_and_727_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_182_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_730_nl = CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_731_nl = CONVOLUTION_LOOP_for_for_for_if_and_549_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_182_nl , CONVOLUTION_LOOP_for_for_for_and_730_nl
      , CONVOLUTION_LOOP_for_for_for_and_731_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_183_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_734_nl = CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_735_nl = CONVOLUTION_LOOP_for_for_for_if_and_551_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_183_nl , CONVOLUTION_LOOP_for_for_for_and_734_nl
      , CONVOLUTION_LOOP_for_for_for_and_735_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_184_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_738_nl = CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_739_nl = CONVOLUTION_LOOP_for_for_for_if_and_553_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_184_nl , CONVOLUTION_LOOP_for_for_for_and_738_nl
      , CONVOLUTION_LOOP_for_for_for_and_739_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_185_nl = (~(CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_742_nl = CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_743_nl = CONVOLUTION_LOOP_for_for_for_if_and_555_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_185_nl , CONVOLUTION_LOOP_for_for_for_and_742_nl
      , CONVOLUTION_LOOP_for_for_for_and_743_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_186_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_746_nl = CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_747_nl = CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_186_nl , CONVOLUTION_LOOP_for_for_for_and_746_nl
      , CONVOLUTION_LOOP_for_for_for_and_747_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_187_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_750_nl = CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_751_nl = CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_187_nl , CONVOLUTION_LOOP_for_for_for_and_750_nl
      , CONVOLUTION_LOOP_for_for_for_and_751_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_188_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_754_nl = CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_755_nl = CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_188_nl , CONVOLUTION_LOOP_for_for_for_and_754_nl
      , CONVOLUTION_LOOP_for_for_for_and_755_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_189_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_758_nl = CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_759_nl = CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_189_nl , CONVOLUTION_LOOP_for_for_for_and_758_nl
      , CONVOLUTION_LOOP_for_for_for_and_759_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_190_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_762_nl = CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_763_nl = CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_190_nl , CONVOLUTION_LOOP_for_for_for_and_762_nl
      , CONVOLUTION_LOOP_for_for_for_and_763_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_191_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_766_nl = CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_767_nl = CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_191_nl , CONVOLUTION_LOOP_for_for_for_and_766_nl
      , CONVOLUTION_LOOP_for_for_for_and_767_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_192_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_770_nl = CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_771_nl = CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_192_nl , CONVOLUTION_LOOP_for_for_for_and_770_nl
      , CONVOLUTION_LOOP_for_for_for_and_771_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_193_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_774_nl = CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_775_nl = CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_193_nl , CONVOLUTION_LOOP_for_for_for_and_774_nl
      , CONVOLUTION_LOOP_for_for_for_and_775_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_194_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_778_nl = CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_779_nl = CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_194_nl , CONVOLUTION_LOOP_for_for_for_and_778_nl
      , CONVOLUTION_LOOP_for_for_for_and_779_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_195_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_782_nl = CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_783_nl = CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_195_nl , CONVOLUTION_LOOP_for_for_for_and_782_nl
      , CONVOLUTION_LOOP_for_for_for_and_783_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_196_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_786_nl = CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_787_nl = CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_196_nl , CONVOLUTION_LOOP_for_for_for_and_786_nl
      , CONVOLUTION_LOOP_for_for_for_and_787_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_197_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_790_nl = CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_791_nl = CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_197_nl , CONVOLUTION_LOOP_for_for_for_and_790_nl
      , CONVOLUTION_LOOP_for_for_for_and_791_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_198_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_794_nl = CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_795_nl = CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_198_nl , CONVOLUTION_LOOP_for_for_for_and_794_nl
      , CONVOLUTION_LOOP_for_for_for_and_795_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_199_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_798_nl = CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_799_nl = CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_199_nl , CONVOLUTION_LOOP_for_for_for_and_798_nl
      , CONVOLUTION_LOOP_for_for_for_and_799_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_200_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_802_nl = CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_803_nl = CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_200_nl , CONVOLUTION_LOOP_for_for_for_and_802_nl
      , CONVOLUTION_LOOP_for_for_for_and_803_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_201_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_806_nl = CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_807_nl = CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_201_nl , CONVOLUTION_LOOP_for_for_for_and_806_nl
      , CONVOLUTION_LOOP_for_for_for_and_807_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_202_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_810_nl = CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_811_nl = CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_202_nl , CONVOLUTION_LOOP_for_for_for_and_810_nl
      , CONVOLUTION_LOOP_for_for_for_and_811_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_203_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_814_nl = CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_815_nl = CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_203_nl , CONVOLUTION_LOOP_for_for_for_and_814_nl
      , CONVOLUTION_LOOP_for_for_for_and_815_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_204_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_818_nl = CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_819_nl = CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_204_nl , CONVOLUTION_LOOP_for_for_for_and_818_nl
      , CONVOLUTION_LOOP_for_for_for_and_819_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_205_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_822_nl = CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_823_nl = CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_205_nl , CONVOLUTION_LOOP_for_for_for_and_822_nl
      , CONVOLUTION_LOOP_for_for_for_and_823_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_206_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_826_nl = CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_827_nl = CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_206_nl , CONVOLUTION_LOOP_for_for_for_and_826_nl
      , CONVOLUTION_LOOP_for_for_for_and_827_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_207_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_830_nl = CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_831_nl = CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_207_nl , CONVOLUTION_LOOP_for_for_for_and_830_nl
      , CONVOLUTION_LOOP_for_for_for_and_831_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_208_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_834_nl = CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_835_nl = CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_208_nl , CONVOLUTION_LOOP_for_for_for_and_834_nl
      , CONVOLUTION_LOOP_for_for_for_and_835_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_209_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_838_nl = CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_839_nl = CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_209_nl , CONVOLUTION_LOOP_for_for_for_and_838_nl
      , CONVOLUTION_LOOP_for_for_for_and_839_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_210_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_842_nl = CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_843_nl = CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_210_nl , CONVOLUTION_LOOP_for_for_for_and_842_nl
      , CONVOLUTION_LOOP_for_for_for_and_843_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_211_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_846_nl = CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_847_nl = CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_211_nl , CONVOLUTION_LOOP_for_for_for_and_846_nl
      , CONVOLUTION_LOOP_for_for_for_and_847_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_212_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_850_nl = CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_851_nl = CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_212_nl , CONVOLUTION_LOOP_for_for_for_and_850_nl
      , CONVOLUTION_LOOP_for_for_for_and_851_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_213_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_854_nl = CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_855_nl = CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_213_nl , CONVOLUTION_LOOP_for_for_for_and_854_nl
      , CONVOLUTION_LOOP_for_for_for_and_855_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_214_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_858_nl = CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_859_nl = CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_214_nl , CONVOLUTION_LOOP_for_for_for_and_858_nl
      , CONVOLUTION_LOOP_for_for_for_and_859_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_215_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_862_nl = CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_863_nl = CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_215_nl , CONVOLUTION_LOOP_for_for_for_and_862_nl
      , CONVOLUTION_LOOP_for_for_for_and_863_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_216_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_866_nl = CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_867_nl = CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_216_nl , CONVOLUTION_LOOP_for_for_for_and_866_nl
      , CONVOLUTION_LOOP_for_for_for_and_867_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_217_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_870_nl = CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_871_nl = CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_217_nl , CONVOLUTION_LOOP_for_for_for_and_870_nl
      , CONVOLUTION_LOOP_for_for_for_and_871_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_218_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_874_nl = CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_875_nl = CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_218_nl , CONVOLUTION_LOOP_for_for_for_and_874_nl
      , CONVOLUTION_LOOP_for_for_for_and_875_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_219_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_878_nl = CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_879_nl = CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_219_nl , CONVOLUTION_LOOP_for_for_for_and_878_nl
      , CONVOLUTION_LOOP_for_for_for_and_879_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_220_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_882_nl = CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_883_nl = CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_220_nl , CONVOLUTION_LOOP_for_for_for_and_882_nl
      , CONVOLUTION_LOOP_for_for_for_and_883_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_221_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_886_nl = CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_887_nl = CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_221_nl , CONVOLUTION_LOOP_for_for_for_and_886_nl
      , CONVOLUTION_LOOP_for_for_for_and_887_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_222_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_890_nl = CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_891_nl = CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_222_nl , CONVOLUTION_LOOP_for_for_for_and_890_nl
      , CONVOLUTION_LOOP_for_for_for_and_891_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_223_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_894_nl = CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_895_nl = CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_223_nl , CONVOLUTION_LOOP_for_for_for_and_894_nl
      , CONVOLUTION_LOOP_for_for_for_and_895_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_224_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_898_nl = CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_899_nl = CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_224_nl , CONVOLUTION_LOOP_for_for_for_and_898_nl
      , CONVOLUTION_LOOP_for_for_for_and_899_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_225_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_902_nl = CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_903_nl = CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_225_nl , CONVOLUTION_LOOP_for_for_for_and_902_nl
      , CONVOLUTION_LOOP_for_for_for_and_903_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_226_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_906_nl = CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_907_nl = CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_226_nl , CONVOLUTION_LOOP_for_for_for_and_906_nl
      , CONVOLUTION_LOOP_for_for_for_and_907_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_227_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_910_nl = CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_911_nl = CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_227_nl , CONVOLUTION_LOOP_for_for_for_and_910_nl
      , CONVOLUTION_LOOP_for_for_for_and_911_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_228_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_914_nl = CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_915_nl = CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_228_nl , CONVOLUTION_LOOP_for_for_for_and_914_nl
      , CONVOLUTION_LOOP_for_for_for_and_915_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_229_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_918_nl = CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_919_nl = CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_229_nl , CONVOLUTION_LOOP_for_for_for_and_918_nl
      , CONVOLUTION_LOOP_for_for_for_and_919_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_230_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_922_nl = CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_923_nl = CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_230_nl , CONVOLUTION_LOOP_for_for_for_and_922_nl
      , CONVOLUTION_LOOP_for_for_for_and_923_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_231_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_926_nl = CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_927_nl = CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_231_nl , CONVOLUTION_LOOP_for_for_for_and_926_nl
      , CONVOLUTION_LOOP_for_for_for_and_927_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_232_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_930_nl = CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_931_nl = CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_232_nl , CONVOLUTION_LOOP_for_for_for_and_930_nl
      , CONVOLUTION_LOOP_for_for_for_and_931_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_233_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_934_nl = CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_935_nl = CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_233_nl , CONVOLUTION_LOOP_for_for_for_and_934_nl
      , CONVOLUTION_LOOP_for_for_for_and_935_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_234_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_938_nl = CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_939_nl = CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_234_nl , CONVOLUTION_LOOP_for_for_for_and_938_nl
      , CONVOLUTION_LOOP_for_for_for_and_939_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_235_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_942_nl = CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_943_nl = CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_235_nl , CONVOLUTION_LOOP_for_for_for_and_942_nl
      , CONVOLUTION_LOOP_for_for_for_and_943_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_236_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_946_nl = CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_947_nl = CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_236_nl , CONVOLUTION_LOOP_for_for_for_and_946_nl
      , CONVOLUTION_LOOP_for_for_for_and_947_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_237_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_950_nl = CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_951_nl = CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_237_nl , CONVOLUTION_LOOP_for_for_for_and_950_nl
      , CONVOLUTION_LOOP_for_for_for_and_951_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_238_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_954_nl = CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_955_nl = CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_238_nl , CONVOLUTION_LOOP_for_for_for_and_954_nl
      , CONVOLUTION_LOOP_for_for_for_and_955_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_239_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_958_nl = CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_959_nl = CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_239_nl , CONVOLUTION_LOOP_for_for_for_and_958_nl
      , CONVOLUTION_LOOP_for_for_for_and_959_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_240_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_962_nl = CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_963_nl = CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_240_nl , CONVOLUTION_LOOP_for_for_for_and_962_nl
      , CONVOLUTION_LOOP_for_for_for_and_963_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_241_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_966_nl = CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_967_nl = CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_241_nl , CONVOLUTION_LOOP_for_for_for_and_966_nl
      , CONVOLUTION_LOOP_for_for_for_and_967_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_242_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_970_nl = CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_971_nl = CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_242_nl , CONVOLUTION_LOOP_for_for_for_and_970_nl
      , CONVOLUTION_LOOP_for_for_for_and_971_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_243_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_974_nl = CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_975_nl = CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_243_nl , CONVOLUTION_LOOP_for_for_for_and_974_nl
      , CONVOLUTION_LOOP_for_for_for_and_975_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_244_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_978_nl = CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_979_nl = CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_244_nl , CONVOLUTION_LOOP_for_for_for_and_978_nl
      , CONVOLUTION_LOOP_for_for_for_and_979_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_245_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_982_nl = CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_983_nl = CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_245_nl , CONVOLUTION_LOOP_for_for_for_and_982_nl
      , CONVOLUTION_LOOP_for_for_for_and_983_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_246_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_986_nl = CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_987_nl = CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_246_nl , CONVOLUTION_LOOP_for_for_for_and_986_nl
      , CONVOLUTION_LOOP_for_for_for_and_987_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_247_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_990_nl = CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_991_nl = CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_247_nl , CONVOLUTION_LOOP_for_for_for_and_990_nl
      , CONVOLUTION_LOOP_for_for_for_and_991_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_248_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_994_nl = CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_995_nl = CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_248_nl , CONVOLUTION_LOOP_for_for_for_and_994_nl
      , CONVOLUTION_LOOP_for_for_for_and_995_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_249_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_998_nl = CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_999_nl = CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_249_nl , CONVOLUTION_LOOP_for_for_for_and_998_nl
      , CONVOLUTION_LOOP_for_for_for_and_999_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_250_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1002_nl = CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1003_nl = CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_250_nl , CONVOLUTION_LOOP_for_for_for_and_1002_nl
      , CONVOLUTION_LOOP_for_for_for_and_1003_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_251_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1006_nl = CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1007_nl = CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_251_nl , CONVOLUTION_LOOP_for_for_for_and_1006_nl
      , CONVOLUTION_LOOP_for_for_for_and_1007_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_252_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1010_nl = CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1011_nl = CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_252_nl , CONVOLUTION_LOOP_for_for_for_and_1010_nl
      , CONVOLUTION_LOOP_for_for_for_and_1011_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_253_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1014_nl = CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1015_nl = CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_253_nl , CONVOLUTION_LOOP_for_for_for_and_1014_nl
      , CONVOLUTION_LOOP_for_for_for_and_1015_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_254_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1018_nl = CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1019_nl = CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_254_nl , CONVOLUTION_LOOP_for_for_for_and_1018_nl
      , CONVOLUTION_LOOP_for_for_for_and_1019_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_255_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1022_nl = CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1023_nl = CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_255_nl , CONVOLUTION_LOOP_for_for_for_and_1022_nl
      , CONVOLUTION_LOOP_for_for_for_and_1023_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_256_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1026_nl = CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1027_nl = CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_256_nl , CONVOLUTION_LOOP_for_for_for_and_1026_nl
      , CONVOLUTION_LOOP_for_for_for_and_1027_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_257_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1030_nl = CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1031_nl = CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_257_nl , CONVOLUTION_LOOP_for_for_for_and_1030_nl
      , CONVOLUTION_LOOP_for_for_for_and_1031_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_258_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1034_nl = CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1035_nl = CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_258_nl , CONVOLUTION_LOOP_for_for_for_and_1034_nl
      , CONVOLUTION_LOOP_for_for_for_and_1035_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_259_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1038_nl = CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1039_nl = CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_259_nl , CONVOLUTION_LOOP_for_for_for_and_1038_nl
      , CONVOLUTION_LOOP_for_for_for_and_1039_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_260_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1042_nl = CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1043_nl = CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_260_nl , CONVOLUTION_LOOP_for_for_for_and_1042_nl
      , CONVOLUTION_LOOP_for_for_for_and_1043_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_261_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1046_nl = CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1047_nl = CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_261_nl , CONVOLUTION_LOOP_for_for_for_and_1046_nl
      , CONVOLUTION_LOOP_for_for_for_and_1047_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_262_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1050_nl = CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1051_nl = CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_262_nl , CONVOLUTION_LOOP_for_for_for_and_1050_nl
      , CONVOLUTION_LOOP_for_for_for_and_1051_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_263_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1054_nl = CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1055_nl = CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_263_nl , CONVOLUTION_LOOP_for_for_for_and_1054_nl
      , CONVOLUTION_LOOP_for_for_for_and_1055_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_264_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1058_nl = CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1059_nl = CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_264_nl , CONVOLUTION_LOOP_for_for_for_and_1058_nl
      , CONVOLUTION_LOOP_for_for_for_and_1059_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_265_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1062_nl = CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1063_nl = CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_265_nl , CONVOLUTION_LOOP_for_for_for_and_1062_nl
      , CONVOLUTION_LOOP_for_for_for_and_1063_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_266_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1066_nl = CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1067_nl = CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_266_nl , CONVOLUTION_LOOP_for_for_for_and_1066_nl
      , CONVOLUTION_LOOP_for_for_for_and_1067_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_267_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1070_nl = CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1071_nl = CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_267_nl , CONVOLUTION_LOOP_for_for_for_and_1070_nl
      , CONVOLUTION_LOOP_for_for_for_and_1071_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_268_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1074_nl = CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1075_nl = CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_268_nl , CONVOLUTION_LOOP_for_for_for_and_1074_nl
      , CONVOLUTION_LOOP_for_for_for_and_1075_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_269_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1078_nl = CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1079_nl = CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_269_nl , CONVOLUTION_LOOP_for_for_for_and_1078_nl
      , CONVOLUTION_LOOP_for_for_for_and_1079_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_270_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1082_nl = CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1083_nl = CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_270_nl , CONVOLUTION_LOOP_for_for_for_and_1082_nl
      , CONVOLUTION_LOOP_for_for_for_and_1083_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_271_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1086_nl = CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1087_nl = CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_271_nl , CONVOLUTION_LOOP_for_for_for_and_1086_nl
      , CONVOLUTION_LOOP_for_for_for_and_1087_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_272_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1090_nl = CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1091_nl = CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_272_nl , CONVOLUTION_LOOP_for_for_for_and_1090_nl
      , CONVOLUTION_LOOP_for_for_for_and_1091_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_273_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1094_nl = CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1095_nl = CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_273_nl , CONVOLUTION_LOOP_for_for_for_and_1094_nl
      , CONVOLUTION_LOOP_for_for_for_and_1095_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_274_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1098_nl = CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1099_nl = CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_274_nl , CONVOLUTION_LOOP_for_for_for_and_1098_nl
      , CONVOLUTION_LOOP_for_for_for_and_1099_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_275_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1102_nl = CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1103_nl = CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_275_nl , CONVOLUTION_LOOP_for_for_for_and_1102_nl
      , CONVOLUTION_LOOP_for_for_for_and_1103_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_276_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1106_nl = CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1107_nl = CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_276_nl , CONVOLUTION_LOOP_for_for_for_and_1106_nl
      , CONVOLUTION_LOOP_for_for_for_and_1107_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_277_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1110_nl = CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1111_nl = CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_277_nl , CONVOLUTION_LOOP_for_for_for_and_1110_nl
      , CONVOLUTION_LOOP_for_for_for_and_1111_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_278_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1114_nl = CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1115_nl = CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_278_nl , CONVOLUTION_LOOP_for_for_for_and_1114_nl
      , CONVOLUTION_LOOP_for_for_for_and_1115_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_279_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1118_nl = CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1119_nl = CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_279_nl , CONVOLUTION_LOOP_for_for_for_and_1118_nl
      , CONVOLUTION_LOOP_for_for_for_and_1119_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_280_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1122_nl = CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1123_nl = CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_280_nl , CONVOLUTION_LOOP_for_for_for_and_1122_nl
      , CONVOLUTION_LOOP_for_for_for_and_1123_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_281_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1126_nl = CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1127_nl = CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_281_nl , CONVOLUTION_LOOP_for_for_for_and_1126_nl
      , CONVOLUTION_LOOP_for_for_for_and_1127_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_282_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1130_nl = CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1131_nl = CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_282_nl , CONVOLUTION_LOOP_for_for_for_and_1130_nl
      , CONVOLUTION_LOOP_for_for_for_and_1131_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_283_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1134_nl = CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1135_nl = CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_283_nl , CONVOLUTION_LOOP_for_for_for_and_1134_nl
      , CONVOLUTION_LOOP_for_for_for_and_1135_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_284_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1138_nl = CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1139_nl = CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_284_nl , CONVOLUTION_LOOP_for_for_for_and_1138_nl
      , CONVOLUTION_LOOP_for_for_for_and_1139_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_285_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1142_nl = CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1143_nl = CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_285_nl , CONVOLUTION_LOOP_for_for_for_and_1142_nl
      , CONVOLUTION_LOOP_for_for_for_and_1143_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_286_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1146_nl = CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1147_nl = CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_286_nl , CONVOLUTION_LOOP_for_for_for_and_1146_nl
      , CONVOLUTION_LOOP_for_for_for_and_1147_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_287_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1150_nl = CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1151_nl = CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_287_nl , CONVOLUTION_LOOP_for_for_for_and_1150_nl
      , CONVOLUTION_LOOP_for_for_for_and_1151_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_288_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1154_nl = CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1155_nl = CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_288_nl , CONVOLUTION_LOOP_for_for_for_and_1154_nl
      , CONVOLUTION_LOOP_for_for_for_and_1155_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_289_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1158_nl = CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1159_nl = CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_289_nl , CONVOLUTION_LOOP_for_for_for_and_1158_nl
      , CONVOLUTION_LOOP_for_for_for_and_1159_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_290_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1162_nl = CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1163_nl = CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_290_nl , CONVOLUTION_LOOP_for_for_for_and_1162_nl
      , CONVOLUTION_LOOP_for_for_for_and_1163_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_291_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1166_nl = CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1167_nl = CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_291_nl , CONVOLUTION_LOOP_for_for_for_and_1166_nl
      , CONVOLUTION_LOOP_for_for_for_and_1167_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_292_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1170_nl = CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1171_nl = CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_292_nl , CONVOLUTION_LOOP_for_for_for_and_1170_nl
      , CONVOLUTION_LOOP_for_for_for_and_1171_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_293_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1174_nl = CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1175_nl = CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_293_nl , CONVOLUTION_LOOP_for_for_for_and_1174_nl
      , CONVOLUTION_LOOP_for_for_for_and_1175_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_294_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1178_nl = CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1179_nl = CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_294_nl , CONVOLUTION_LOOP_for_for_for_and_1178_nl
      , CONVOLUTION_LOOP_for_for_for_and_1179_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_295_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1182_nl = CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1183_nl = CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_295_nl , CONVOLUTION_LOOP_for_for_for_and_1182_nl
      , CONVOLUTION_LOOP_for_for_for_and_1183_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_296_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1186_nl = CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1187_nl = CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_296_nl , CONVOLUTION_LOOP_for_for_for_and_1186_nl
      , CONVOLUTION_LOOP_for_for_for_and_1187_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_297_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1190_nl = CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1191_nl = CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_297_nl , CONVOLUTION_LOOP_for_for_for_and_1190_nl
      , CONVOLUTION_LOOP_for_for_for_and_1191_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_298_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1194_nl = CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1195_nl = CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_298_nl , CONVOLUTION_LOOP_for_for_for_and_1194_nl
      , CONVOLUTION_LOOP_for_for_for_and_1195_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_299_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1198_nl = CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1199_nl = CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_299_nl , CONVOLUTION_LOOP_for_for_for_and_1198_nl
      , CONVOLUTION_LOOP_for_for_for_and_1199_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_300_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1202_nl = CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1203_nl = CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_300_nl , CONVOLUTION_LOOP_for_for_for_and_1202_nl
      , CONVOLUTION_LOOP_for_for_for_and_1203_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_301_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1206_nl = CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1207_nl = CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_301_nl , CONVOLUTION_LOOP_for_for_for_and_1206_nl
      , CONVOLUTION_LOOP_for_for_for_and_1207_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_302_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1210_nl = CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1211_nl = CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_302_nl , CONVOLUTION_LOOP_for_for_for_and_1210_nl
      , CONVOLUTION_LOOP_for_for_for_and_1211_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_303_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1214_nl = CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1215_nl = CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_303_nl , CONVOLUTION_LOOP_for_for_for_and_1214_nl
      , CONVOLUTION_LOOP_for_for_for_and_1215_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_304_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1218_nl = CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1219_nl = CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_304_nl , CONVOLUTION_LOOP_for_for_for_and_1218_nl
      , CONVOLUTION_LOOP_for_for_for_and_1219_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_305_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1222_nl = CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1223_nl = CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_305_nl , CONVOLUTION_LOOP_for_for_for_and_1222_nl
      , CONVOLUTION_LOOP_for_for_for_and_1223_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_306_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1226_nl = CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1227_nl = CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_306_nl , CONVOLUTION_LOOP_for_for_for_and_1226_nl
      , CONVOLUTION_LOOP_for_for_for_and_1227_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_307_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1230_nl = CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1231_nl = CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_307_nl , CONVOLUTION_LOOP_for_for_for_and_1230_nl
      , CONVOLUTION_LOOP_for_for_for_and_1231_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_308_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1234_nl = CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1235_nl = CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_308_nl , CONVOLUTION_LOOP_for_for_for_and_1234_nl
      , CONVOLUTION_LOOP_for_for_for_and_1235_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_309_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1238_nl = CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1239_nl = CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_309_nl , CONVOLUTION_LOOP_for_for_for_and_1238_nl
      , CONVOLUTION_LOOP_for_for_for_and_1239_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_310_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1242_nl = CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1243_nl = CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_310_nl , CONVOLUTION_LOOP_for_for_for_and_1242_nl
      , CONVOLUTION_LOOP_for_for_for_and_1243_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_311_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1246_nl = CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1247_nl = CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_311_nl , CONVOLUTION_LOOP_for_for_for_and_1246_nl
      , CONVOLUTION_LOOP_for_for_for_and_1247_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_312_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1250_nl = CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1251_nl = CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_312_nl , CONVOLUTION_LOOP_for_for_for_and_1250_nl
      , CONVOLUTION_LOOP_for_for_for_and_1251_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_313_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1254_nl = CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1255_nl = CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_313_nl , CONVOLUTION_LOOP_for_for_for_and_1254_nl
      , CONVOLUTION_LOOP_for_for_for_and_1255_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_314_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1258_nl = CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1259_nl = CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_314_nl , CONVOLUTION_LOOP_for_for_for_and_1258_nl
      , CONVOLUTION_LOOP_for_for_for_and_1259_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_315_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1262_nl = CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1263_nl = CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_315_nl , CONVOLUTION_LOOP_for_for_for_and_1262_nl
      , CONVOLUTION_LOOP_for_for_for_and_1263_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_316_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1266_nl = CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1267_nl = CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_316_nl , CONVOLUTION_LOOP_for_for_for_and_1266_nl
      , CONVOLUTION_LOOP_for_for_for_and_1267_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_317_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1270_nl = CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1271_nl = CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_317_nl , CONVOLUTION_LOOP_for_for_for_and_1270_nl
      , CONVOLUTION_LOOP_for_for_for_and_1271_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_318_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1274_nl = CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1275_nl = CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_318_nl , CONVOLUTION_LOOP_for_for_for_and_1274_nl
      , CONVOLUTION_LOOP_for_for_for_and_1275_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_319_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1278_nl = CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1279_nl = CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_319_nl , CONVOLUTION_LOOP_for_for_for_and_1278_nl
      , CONVOLUTION_LOOP_for_for_for_and_1279_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_320_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1282_nl = CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1283_nl = CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_320_nl , CONVOLUTION_LOOP_for_for_for_and_1282_nl
      , CONVOLUTION_LOOP_for_for_for_and_1283_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_321_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1286_nl = CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1287_nl = CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_321_nl , CONVOLUTION_LOOP_for_for_for_and_1286_nl
      , CONVOLUTION_LOOP_for_for_for_and_1287_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_322_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1290_nl = CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1291_nl = CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_322_nl , CONVOLUTION_LOOP_for_for_for_and_1290_nl
      , CONVOLUTION_LOOP_for_for_for_and_1291_nl});
  assign CONVOLUTION_LOOP_for_for_for_or_323_nl = (~(CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1294_nl = CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_and_1295_nl = CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1_dfm_2 = MUX1HOT_v_55_3_2(COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1,
      CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_55_1_sva_1,
      {CONVOLUTION_LOOP_for_for_for_or_323_nl , CONVOLUTION_LOOP_for_for_for_and_1294_nl
      , CONVOLUTION_LOOP_for_for_for_and_1295_nl});
  assign nl_operator_8_false_3_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_135_128_mx0)
      + 9'b111111111;
  assign operator_8_false_3_acc_tmp = nl_operator_8_false_3_acc_tmp[8:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1
      + 5'b00001;
  assign CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2[4:0];
  assign nl_operator_8_false_4_acc_tmp = conv_u2s_8_9(n_h_out_lpi_1_dfm_2) + 9'b111111111;
  assign operator_8_false_4_acc_tmp = nl_operator_8_false_4_acc_tmp[8:0];
  assign if_mux_6_nl = MUX_v_8_2_2(if_acc_4_cse_1, (else_acc_2_psp_sva_1[8:1]), or_314_cse);
  assign operator_42_true_1_and_1_nl = (else_acc_2_psp_sva_1[10]) & (else_acc_2_psp_sva_1[0]);
  assign if_mux_7_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[47:40]), ({7'b0000000
      , operator_42_true_1_and_1_nl}), or_314_cse);
  assign nl_acc_4_nl = ({if_mux_6_nl , 1'b1}) + ({if_mux_7_nl , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[8:0];
  assign n_h_out_lpi_1_dfm_2 = MUX_v_8_2_2(n_h_out_lpi_1_dfm_1, (readslicef_9_8_1(acc_4_nl)),
      COMPUTE_LOOP_or_2_cse);
  assign conf_info_crt_lpi_1_dfm_135_128_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_135_128,
      (conf_info_rsci_idat_mxwt[39:32]), exitL_exit_COMPUTE_LOOP_sva);
  assign CONVOLUTION_LOOP_for_for_for_unequal_tmp_1 = (CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0!=5'b00000);
  assign exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0 = ~(operator_8_false_5_acc_itm_3_1
      & ((~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp))
      | (operator_8_false_1_acc_tmp[8])));
  assign nl_operator_8_false_5_acc_nl = ({1'b1 , CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2})
      + 4'b0001;
  assign operator_8_false_5_acc_nl = nl_operator_8_false_5_acc_nl[3:0];
  assign operator_8_false_5_acc_itm_3_1 = readslicef_4_1_3(operator_8_false_5_acc_nl);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2 = CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_1
      + 3'b001;
  assign CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2[2:0];
  assign CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp = CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_1
      == (operator_8_false_1_acc_tmp[2:0]);
  assign nl_operator_8_false_1_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_103_96_mx0)
      + 9'b111111111;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[8:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp = ~((operator_8_false_1_acc_tmp[7:3]!=5'b00000));
  assign nl_operator_8_false_6_acc_nl = ({1'b1 , CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2})
      + 4'b0001;
  assign operator_8_false_6_acc_nl = nl_operator_8_false_6_acc_nl[3:0];
  assign operator_8_false_6_acc_itm_3_1 = readslicef_4_1_3(operator_8_false_6_acc_nl);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2 = CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_1
      + 3'b001;
  assign CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2[2:0];
  assign CONVOLUTION_LOOP_for_for_for_for_mux_974_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0,
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1, and_tmp_13);
  assign exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_4 = CONVOLUTION_LOOP_for_for_for_for_mux_974_nl
      & exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_1_dfm_1;
  assign exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_1_dfm_1 = ~(operator_8_false_6_acc_itm_3_1
      & ((~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp))
      | (operator_8_false_1_acc_tmp[8])));
  assign CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp = CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_1
      == (operator_8_false_1_acc_tmp[2:0]);
  assign conf_info_crt_lpi_1_dfm_103_96_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_103_96,
      (conf_info_rsci_idat_mxwt[31:24]), exitL_exit_COMPUTE_LOOP_sva);
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_nl = (CONVOLUTION_LOOP_for_for_for_for_for_mul_1_sdt_sva_1[15])
      & ((CONVOLUTION_LOOP_for_for_for_for_for_mul_1_sdt_sva_1[14:0]!=15'b000000000000000)
      | (CONVOLUTION_LOOP_for_for_for_for_for_acc_5_psp_sva_1[0]));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1 = CONVOLUTION_LOOP_for_for_for_for_for_acc_5_psp_sva_1
      + conv_u2s_1_58(CONVOLUTION_LOOP_for_for_for_for_for_and_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1[57:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1[57:56]==2'b10);
  assign CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_for_for_acc_2_psp_sva_1[57:56]!=2'b01));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_5_psp_sva_1 = conv_s2u_57_58({CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
      , CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
      , CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1})
      + conv_s2u_48_58(CONVOLUTION_LOOP_for_for_for_for_for_mul_1_sdt_sva_1[63:16]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_5_psp_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_5_psp_sva_1[57:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_nl = ({CONVOLUTION_LOOP_for_for_for_for_for_x_tmp_2_0_lpi_1_dfm_1
      , CONVOLUTION_LOOP_for_for_for_for_for_x_tmp_2_0_lpi_1_dfm_1}) + (CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1_dfm_mx0[6:1]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_nl[5:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_7_nl = MUX_v_32_126_2((COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[31:0]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[63:32]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[95:64]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[127:96]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[159:128]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[191:160]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[223:192]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[255:224]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[287:256]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[319:288]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[351:320]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[383:352]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[415:384]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[447:416]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[479:448]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[511:480]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[543:512]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[575:544]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[607:576]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[639:608]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[671:640]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[703:672]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[735:704]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[767:736]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[799:768]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[831:800]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[863:832]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[895:864]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[927:896]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[959:928]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[991:960]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1023:992]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1055:1024]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1087:1056]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1119:1088]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1151:1120]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1183:1152]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1215:1184]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1247:1216]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1279:1248]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1311:1280]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1343:1312]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1375:1344]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1407:1376]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1439:1408]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1471:1440]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1503:1472]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1535:1504]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1567:1536]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1599:1568]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1631:1600]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1663:1632]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1695:1664]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1727:1696]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1759:1728]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1791:1760]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1823:1792]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1855:1824]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1887:1856]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1919:1888]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1951:1920]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[1983:1952]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2015:1984]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2047:2016]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2079:2048]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2111:2080]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2143:2112]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2175:2144]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2207:2176]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2239:2208]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2271:2240]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2303:2272]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2335:2304]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2367:2336]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2399:2368]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2431:2400]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2463:2432]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2495:2464]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2527:2496]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2559:2528]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2591:2560]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2623:2592]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2655:2624]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2687:2656]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2719:2688]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2751:2720]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2783:2752]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2815:2784]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2847:2816]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2879:2848]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2911:2880]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2943:2912]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[2975:2944]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3007:2976]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3039:3008]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3071:3040]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3103:3072]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3135:3104]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3167:3136]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3199:3168]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3231:3200]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3263:3232]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3295:3264]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3327:3296]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3359:3328]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3391:3360]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3423:3392]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3455:3424]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3487:3456]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3519:3488]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3551:3520]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3583:3552]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3615:3584]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3647:3616]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3679:3648]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3711:3680]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3743:3712]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3775:3744]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3807:3776]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3839:3808]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3871:3840]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3903:3872]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3935:3904]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3967:3936]), (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[3999:3968]),
      (COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0[4031:4000]), {CONVOLUTION_LOOP_for_for_for_for_for_acc_nl
      , (CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1_dfm_mx0[0])});
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_index_f_mul_nl = CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_1
      * (conf_info_crt_lpi_1_dfm_103_96_mx0[5:0]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_index_f_mul_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_index_f_mul_nl[5:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_index_f_acc_nl = CONVOLUTION_LOOP_for_for_for_for_for_index_f_mul_nl
      + conv_u2u_3_6(CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_1);
  assign CONVOLUTION_LOOP_for_for_for_for_for_index_f_acc_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_index_f_acc_nl[5:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_8_nl = MUX_v_32_49_2((COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[31:0]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[63:32]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[95:64]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[127:96]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[159:128]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[191:160]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[223:192]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[255:224]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[287:256]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[319:288]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[351:320]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[383:352]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[415:384]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[447:416]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[479:448]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[511:480]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[543:512]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[575:544]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[607:576]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[639:608]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[671:640]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[703:672]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[735:704]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[767:736]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[799:768]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[831:800]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[863:832]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[895:864]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[927:896]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[959:928]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[991:960]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1023:992]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1055:1024]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1087:1056]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1119:1088]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1151:1120]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1183:1152]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1215:1184]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1247:1216]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1279:1248]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1311:1280]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1343:1312]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1375:1344]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1407:1376]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1439:1408]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1471:1440]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1503:1472]),
      (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1535:1504]), (COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0[1567:1536]),
      CONVOLUTION_LOOP_for_for_for_for_for_index_f_acc_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_1_sdt_sva_1 = conv_s2u_64_64($signed(CONVOLUTION_LOOP_for_for_for_for_for_mux_7_nl)
      * $signed(CONVOLUTION_LOOP_for_for_for_for_for_mux_8_nl));
  assign COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm_mx0 = MUX_v_4032_2_2(COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm,
      buf_linear_rsci_idat_mxwt, exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1);
  assign nl_operator_8_false_1_acc_3_nl = conv_u2u_1_2(operator_8_false_1_acc_imod_2_sva_1[0])
      + conv_u2u_1_2(operator_8_false_1_acc_imod_2_sva_1[1]);
  assign operator_8_false_1_acc_3_nl = nl_operator_8_false_1_acc_3_nl[1:0];
  assign nl_operator_8_false_2_acc_2_nl = conv_u2u_1_3(z_out_2_2_0[2]) + conv_u2u_2_3(z_out_2_2_0[1:0]);
  assign operator_8_false_2_acc_2_nl = nl_operator_8_false_2_acc_2_nl[2:0];
  assign nl_operator_8_false_3_operator_8_false_3_acc_nl = conv_s2u_1_3(z_out_2_2_0[2])
      + z_out_2_2_0;
  assign operator_8_false_3_operator_8_false_3_acc_nl = nl_operator_8_false_3_operator_8_false_3_acc_nl[2:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_and_3_nl
      = (conf_info_crt_lpi_1_dfm_103_96_mx0==8'b00000111);
  assign CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_mux1h_7_nl = MUX1HOT_v_3_3_2(({1'b0
      , operator_8_false_1_acc_3_nl}), operator_8_false_2_acc_2_nl, operator_8_false_3_operator_8_false_3_acc_nl,
      {(~ (conf_info_crt_lpi_1_dfm_103_96_mx0[2])) , (~ (conf_info_crt_lpi_1_dfm_103_96_mx0[1]))
      , CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_and_3_nl});
  assign CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_nand_nl
      = ~((conf_info_crt_lpi_1_dfm_103_96_mx0==8'b00000001));
  assign CONVOLUTION_LOOP_for_for_for_for_for_x_tmp_2_0_lpi_1_dfm_1 = MUX_v_3_2_2(3'b000,
      CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_mux1h_7_nl, CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_CONVOLUTION_LOOP_for_for_for_for_for_switch_lp_nand_nl);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1
      * (conf_info_crt_lpi_1_dfm_7_0_mx0[6:0]);
  assign CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0 = nl_CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0[6:0];
  assign CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1_dfm_mx0 = MUX_v_7_2_2(CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1,
      CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0, exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1);
  assign COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm_mx0 = MUX_v_1568_2_2(COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm,
      plm_kernel_rsci_idat_mxwt, exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1);
  assign exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0 = (exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_4
      & main_stage_v_1) | exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1;
  assign nand_76_cse = ~(main_stage_v_2 & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1
      & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
      & (~ var_output_rsci_bawt));
  assign or_61_cse = (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1) |
      (~ CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1)
      | var_output_rsci_bawt;
  assign or_dcpl_11 = done_rsci_bawt | (~ exit_COMPUTE_LOOP_lpi_1_dfm_3_st_2);
  assign or_dcpl_12 = or_dcpl_11 | (~ main_stage_v_3);
  assign and_dcpl_8 = or_dcpl_12 & or_61_cse;
  assign and_dcpl_13 = (~ var_output_rsci_bawt) & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1;
  assign and_dcpl_14 = (and_dcpl_13 | (~ main_stage_v_2) | (~ exit_COMPUTE_LOOP_lpi_1_dfm_3_st_1))
      & asn_done_rsci_oswt_and_cse;
  assign nand_68_nl = ~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp
      & (~ (operator_8_false_1_acc_tmp[8])) & nand_76_cse);
  assign mux_tmp_27 = MUX_s_1_2_2((~ nand_76_cse), nand_68_nl, operator_8_false_6_acc_itm_3_1);
  assign nand_24_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_42_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8])
      | (~ nand_76_cse))));
  assign mux_tmp_28 = MUX_s_1_2_2(mux_tmp_27, nand_24_nl, operator_8_false_5_acc_itm_3_1);
  assign and_dcpl_25 = (~ mux_tmp_28) & or_dcpl_12 & or_59_cse & or_58_cse & or_57_cse;
  assign and_dcpl_30 = (~ buf_linear_rsci_bawt) & exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1;
  assign and_dcpl_31 = (~ plm_kernel_rsci_bawt) & exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1;
  assign and_dcpl_32 = (~ conf_info_rsci_bawt) & COMPUTE_LOOP_asn_itm_1;
  assign and_tmp_13 = operator_8_false_6_acc_itm_3_1 & or_41_cse;
  assign nand_25_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_42_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8]))));
  assign mux_tmp_29 = MUX_s_1_2_2(and_tmp_13, nand_25_nl, operator_8_false_5_acc_itm_3_1);
  assign and_dcpl_34 = (mux_tmp_29 | and_dcpl_32 | (operator_8_false_3_acc_tmp[8:5]!=4'b0000)
      | and_dcpl_31 | and_dcpl_30 | (~(CONVOLUTION_LOOP_for_if_equal_tmp & main_stage_v_1)))
      & or_dcpl_12 & var_output_rsci_bawt & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1 & main_stage_v_2;
  assign or_dcpl_32 = and_dcpl_31 | and_dcpl_30;
  assign or_dcpl_33 = or_dcpl_32 | (~ main_stage_v_1);
  assign or_dcpl_36 = mux_tmp_28 | and_6_cse | and_dcpl_32;
  assign or_dcpl_38 = and_dcpl_30 | (~ main_stage_v_1);
  assign or_dcpl_42 = (~ nand_76_cse) | and_6_cse;
  assign and_tmp_14 = (done_rsci_bawt | (~ exit_COMPUTE_LOOP_lpi_1_dfm_3_st_2) |
      (~ main_stage_v_3)) & nand_76_cse;
  assign not_tmp_46 = ~(or_57_cse & or_58_cse & and_tmp_14);
  assign nor_32_cse = ~((~ CONVOLUTION_LOOP_for_if_equal_tmp) | (operator_8_false_3_acc_tmp[8:5]!=4'b0000));
  assign and_62_nl = operator_8_false_6_acc_itm_3_1 & or_41_cse & nand_76_cse;
  assign and_60_nl = (nor_42_cse | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)
      | (operator_8_false_1_acc_tmp[8])) & nand_76_cse;
  assign mux_49_nl = MUX_s_1_2_2(nand_76_cse, and_60_nl, CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp);
  assign mux_50_cse = MUX_s_1_2_2(and_62_nl, mux_49_nl, operator_8_false_5_acc_itm_3_1);
  assign mux_51_nl = MUX_s_1_2_2(nand_76_cse, mux_50_cse, or_163_cse);
  assign mux_52_nl = MUX_s_1_2_2(nand_76_cse, mux_51_nl, nand_74_cse);
  assign mux_53_nl = MUX_s_1_2_2(nand_76_cse, mux_52_nl, nand_52_cse);
  assign mux_54_nl = MUX_s_1_2_2(nand_76_cse, mux_53_nl, or_157_cse);
  assign mux_55_nl = MUX_s_1_2_2(nand_76_cse, mux_54_nl, or_155_cse);
  assign and_dcpl_40 = mux_55_nl & or_dcpl_12 & or_58_cse & or_57_cse & conf_info_rsci_bawt
      & COMPUTE_LOOP_asn_itm_1 & main_stage_v_1;
  assign and_tmp_28 = or_57_cse & or_58_cse & or_59_cse & nand_76_cse;
  assign and_143_nl = CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp
      & (~ (operator_8_false_1_acc_tmp[8])) & and_tmp_28;
  assign mux_60_nl = MUX_s_1_2_2(and_tmp_28, and_143_nl, operator_8_false_6_acc_itm_3_1);
  assign and_144_nl = CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_42_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8])
      | (~ and_tmp_28)));
  assign mux_61_nl = MUX_s_1_2_2(mux_60_nl, and_144_nl, operator_8_false_5_acc_itm_3_1);
  assign nand_tmp_20 = ~(nand_74_cse & mux_61_nl);
  assign and_tmp_29 = exitL_exit_COMPUTE_LOOP_sva & nand_76_cse;
  assign mux_66_cse_1 = MUX_s_1_2_2(nand_76_cse, mux_50_cse, nand_74_cse);
  assign mux_96_nl = MUX_s_1_2_2(nand_76_cse, mux_50_cse, nand_74_cse);
  assign mux_67_nl = MUX_s_1_2_2(mux_96_nl, nand_76_cse, or_289_cse);
  assign mux_68_nl = MUX_s_1_2_2(mux_66_cse_1, mux_67_nl, operator_8_false_3_acc_itm_4_1);
  assign and_dcpl_47 = mux_68_nl & or_dcpl_12 & or_59_cse & or_57_cse & plm_kernel_rsci_bawt
      & exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1 & main_stage_v_1;
  assign or_dcpl_51 = and_dcpl_32 | and_dcpl_31;
  assign and_dcpl_54 = mux_66_cse_1 & or_dcpl_12 & or_59_cse & or_58_cse & buf_linear_rsci_bawt
      & exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1 & main_stage_v_1;
  assign mux_78_nl = MUX_s_1_2_2(nand_76_cse, and_tmp_28, main_stage_v_1);
  assign or_dcpl_57 = (~ mux_78_nl) | and_6_cse;
  assign and_dcpl_55 = ~(exit_CONVOLUTION_LOOP_sva_3 | (CONVOLUTION_LOOP_acc_tmp[5]));
  assign and_dcpl_56 = or_289_cse & operator_8_false_3_acc_itm_4_1;
  assign and_dcpl_57 = or_290_cse & operator_8_false_4_acc_itm_4_1;
  assign nand_49_nl = ~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp
      & (~ (operator_8_false_1_acc_tmp[8])) & or_163_cse);
  assign mux_79_nl = MUX_s_1_2_2((~ or_163_cse), nand_49_nl, operator_8_false_6_acc_itm_3_1);
  assign nand_46_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_42_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8])
      | (~ or_163_cse))));
  assign mux_80_nl = MUX_s_1_2_2(mux_79_nl, nand_46_nl, operator_8_false_5_acc_itm_3_1);
  assign or_dcpl_62 = mux_80_nl | and_dcpl_57 | and_dcpl_56;
  assign or_dcpl_63 = or_dcpl_62 | and_dcpl_55;
  assign not_tmp_91 = ~(nand_76_cse & or_163_cse);
  assign or_244_nl = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)
      | (operator_8_false_1_acc_tmp[8]) | not_tmp_91;
  assign mux_81_nl = MUX_s_1_2_2(not_tmp_91, or_244_nl, operator_8_false_6_acc_itm_3_1);
  assign nand_47_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_42_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8])
      | not_tmp_91)));
  assign mux_82_nl = MUX_s_1_2_2(mux_81_nl, nand_47_nl, operator_8_false_5_acc_itm_3_1);
  assign or_dcpl_64 = mux_82_nl | and_6_cse;
  assign or_dcpl_75 = mux_tmp_29 | and_dcpl_57;
  assign or_dcpl_76 = or_dcpl_75 | and_dcpl_56;
  assign and_dcpl_61 = (CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0==5'b00000);
  assign and_dcpl_66 = (~ mux_tmp_27) & or_dcpl_12 & or_59_cse & or_58_cse & or_57_cse
      & main_stage_v_1;
  assign and_dcpl_68 = nand_76_cse & or_dcpl_12;
  assign and_dcpl_71 = and_dcpl_68 & or_59_cse & or_58_cse & or_57_cse;
  assign and_dcpl_73 = and_dcpl_71 & or_41_cse & operator_8_false_6_acc_itm_3_1 &
      main_stage_v_1;
  assign and_dcpl_74 = and_dcpl_71 & main_stage_v_1;
  assign COMPUTE_LOOP_asn_itm_1_mx0c1 = and_dcpl_68 & (~ main_stage_v_1);
  assign main_stage_v_2_mx0c1 = (or_dcpl_51 | or_dcpl_38) & or_dcpl_12 & or_61_cse
      & main_stage_v_2;
  assign CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1
      = mux_50_cse & or_dcpl_12 & or_59_cse & or_58_cse & or_57_cse & main_stage_v_1;
  assign main_stage_v_3_mx0c1 = (and_dcpl_13 | (~ main_stage_v_2)) & or_dcpl_11 &
      main_stage_v_3;
  assign nl_operator_8_false_3_acc_nl = conv_u2s_4_5(CONVOLUTION_LOOP_for_for_i_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_3_acc_nl = nl_operator_8_false_3_acc_nl[4:0];
  assign operator_8_false_3_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_3_acc_nl);
  assign nl_operator_8_false_4_acc_nl = conv_u2s_4_5(CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_4_acc_nl = nl_operator_8_false_4_acc_nl[4:0];
  assign operator_8_false_4_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_4_acc_nl);
  assign or_314_cse = (conf_info_rsci_idat_mxwt[7:0]!=8'b00000001);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_done_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_8 & main_stage_v_2 & exit_COMPUTE_LOOP_lpi_1_dfm_3_st_1)
        | and_dcpl_14) ) begin
      reg_done_rsci_iswt0_cse <= ~ and_dcpl_14;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_var_output_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_25 & (operator_8_false_3_acc_tmp[8:5]==4'b0000)
        & CONVOLUTION_LOOP_for_if_equal_tmp & main_stage_v_1) | and_dcpl_34) ) begin
      reg_var_output_rsci_iswt0_cse <= ~ and_dcpl_34;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      var_output_rsci_idat_31 <= 1'b0;
      var_output_rsci_idat_0 <= 1'b0;
      var_output_rsci_idat_30_1 <= 30'b000000000000000000000000000000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_if_1_and_6_cse ) begin
      var_output_rsci_idat_31 <= ~((~((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_55_1_1[30])
          | CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1);
      var_output_rsci_idat_0 <= ~((~(CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl |
          CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1);
      var_output_rsci_idat_30_1 <= ~(MUX_v_30_2_2(CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl,
          30'b111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1));
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (mux_48_nl | and_dcpl_40) ) begin
      reg_conf_info_rsci_iswt0_cse <= ~ and_dcpl_40;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_kernel_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((mux_63_nl & or_dcpl_12) | and_dcpl_47) ) begin
      reg_plm_kernel_rsci_iswt0_cse <= ~ and_dcpl_47;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_buf_linear_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((mux_73_nl & or_dcpl_12) | and_dcpl_54) ) begin
      reg_buf_linear_rsci_iswt0_cse <= ~ and_dcpl_54;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exitL_exit_COMPUTE_LOOP_sva <= 1'b1;
      n_w_out_lpi_1_dfm_1 <= 8'b00000000;
      n_h_out_lpi_1_dfm_1 <= 8'b00000000;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1 <= 1'b0;
    end
    else if ( COMPUTE_LOOP_and_2_cse ) begin
      exitL_exit_COMPUTE_LOOP_sva <= exit_COMPUTE_LOOP_lpi_1_dfm_3_mx0w0;
      n_w_out_lpi_1_dfm_1 <= n_w_out_lpi_1_dfm_2;
      n_h_out_lpi_1_dfm_1 <= n_h_out_lpi_1_dfm_2;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_1 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_4;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_1 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
          <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
          <= 55'b0000000000000000000000000000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1
          <= 1'b0;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= 1'b0;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1 <= 1'b0;
      exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( and_156_cse ) begin
      main_stage_v_1 <= 1'b1;
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_1 <= MUX_v_3_2_2(3'b000,
          CONVOLUTION_LOOP_for_for_for_for_for_mux_4_nl, CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_not_nl);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
          <= CONVOLUTION_LOOP_for_for_for_acc_56_sva_2 & main_stage_v_1 & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
          <= MUX_v_55_2_2(55'b0000000000000000000000000000000000000000000000000000000,
          CONVOLUTION_LOOP_for_for_for_acc_55_1_sva_2, CONVOLUTION_LOOP_for_for_for_for_not_26_nl);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1
          <= CONVOLUTION_LOOP_for_for_for_acc_0_sva_2 & main_stage_v_1 & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0);
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1 <= exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1;
      exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1 <= exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1 <= 5'b00000;
    end
    else if ( core_wen & (~(((~ exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1)
        & mux_tmp_29) | or_dcpl_57)) ) begin
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1 <= MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2,
          CONVOLUTION_LOOP_for_for_for_not_339_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_crt_lpi_1_dfm_7_0 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_231_224 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_71_64 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_135_128 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_103_96 <= 8'b00000000;
    end
    else if ( core_wen ) begin
      conf_info_crt_lpi_1_dfm_7_0 <= conf_info_crt_lpi_1_dfm_7_0_mx0;
      conf_info_crt_lpi_1_dfm_231_224 <= conf_info_crt_lpi_1_dfm_231_224_mx0;
      conf_info_crt_lpi_1_dfm_71_64 <= conf_info_crt_lpi_1_dfm_71_64_mx0;
      conf_info_crt_lpi_1_dfm_135_128 <= conf_info_crt_lpi_1_dfm_135_128_mx0;
      conf_info_crt_lpi_1_dfm_103_96 <= conf_info_crt_lpi_1_dfm_103_96_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1 <= 5'b00000;
    end
    else if ( core_wen & (~(((~ exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1)
        & or_dcpl_75) | or_dcpl_57)) ) begin
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_1 <= MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_for_i_4_0_sva_2,
          CONVOLUTION_LOOP_for_for_not_14_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_64 | and_dcpl_32 | and_dcpl_57 | and_dcpl_56
        | and_dcpl_55 | and_dcpl_31 | or_dcpl_38)) ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_1 <= or_155_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_LOOP_b_4_0_lpi_1_dfm_1_3_0 <= 4'b0000;
    end
    else if ( core_wen & (~(((~ exitL_exit_COMPUTE_LOOP_sva_mx0) & or_dcpl_63) |
        or_dcpl_57)) ) begin
      COMPUTE_LOOP_b_4_0_lpi_1_dfm_1_3_0 <= MUX_v_4_2_2(4'b0000, (COMPUTE_LOOP_acc_tmp[3:0]),
          COMPUTE_LOOP_not_19_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_64 | or_dcpl_51 | and_dcpl_57 | and_dcpl_56 |
        or_dcpl_38)) ) begin
      exit_CONVOLUTION_LOOP_lpi_1_dfm_1 <= or_157_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_1_4_0 <= 5'b00000;
    end
    else if ( core_wen & (~(((~ exitL_exit_COMPUTE_LOOP_sva_mx0) & or_dcpl_62) |
        or_dcpl_57)) ) begin
      CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_1_4_0 <= MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_CONVOLUTION_LOOP_CONVOLUTION_LOOP_mux_nl,
          COMPUTE_LOOP_COMPUTE_LOOP_COMPUTE_LOOP_COMPUTE_LOOP_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0 <= 5'b00000;
    end
    else if ( core_wen & (~((lfst_exit_CONVOLUTION_LOOP_1_lpi_1_dfm_1 & or_dcpl_76)
        | or_dcpl_57)) ) begin
      CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0 <= MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_mux_nl,
          lfst_exit_CONVOLUTION_LOOP_1_lpi_1_dfm_1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_36 | or_dcpl_32 | and_dcpl_57 | and_dcpl_56 |
        (~ main_stage_v_1))) ) begin
      exit_CONVOLUTION_LOOP_for_sva_2 <= exit_CONVOLUTION_LOOP_for_sva_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1 <= 1'b0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1 <= 55'b0000000000000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm
          <= 1'b0;
    end
    else if ( COMPUTE_LOOP_buf_tmp_acc_data_and_cse ) begin
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_17_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_0_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_16_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_1_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_15_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_2_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_14_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_3_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_13_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_4_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_12_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_5_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_11_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_6_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_10_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_7_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_17_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_8_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_8_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_9_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_9_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_7_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_7_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_10_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_10_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_6_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_6_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_11_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_11_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_5_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_5_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_12_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_12_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_4_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_4_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_13_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_13_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_3_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_3_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_14_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_14_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_2_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_2_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_15_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_15_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_1_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_1_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_16_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_16_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_0_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_9_0_56_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_17_55_1_lpi_1_dfm_2;
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1 <= COMPUTE_LOOP_buf_tmp_acc_data_8_17_56_lpi_1_dfm_1_mx0;
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm
          <= exit_CONVOLUTION_LOOP_for_sva_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(mux_tmp_27 | and_6_cse | and_dcpl_32 | or_dcpl_33)) )
        begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_1 <= 3'b000;
    end
    else if ( core_wen & (~(((~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0)
        & and_tmp_13) | or_dcpl_57)) ) begin
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_1 <= MUX_v_3_2_2(3'b000, CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2,
          CONVOLUTION_LOOP_for_for_for_for_not_22_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1 <= 7'b0000000;
    end
    else if ( core_wen & (CONVOLUTION_LOOP_for_for_for_for_for_and_2_rgt | CONVOLUTION_LOOP_for_for_for_for_for_and_3_rgt
        | and_dcpl_73) ) begin
      CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1 <= MUX1HOT_v_7_3_2(CONVOLUTION_LOOP_for_for_for_y_mul_cse_6_0_lpi_1_dfm,
          CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0, (z_out_5[6:0]), {CONVOLUTION_LOOP_for_for_for_for_for_and_2_rgt
          , CONVOLUTION_LOOP_for_for_for_for_for_and_3_rgt , and_dcpl_73});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_x_lpi_1 <= 8'b00000000;
    end
    else if ( core_wen & (and_dcpl_66 | CONVOLUTION_LOOP_for_for_for_for_for_and_5_rgt)
        ) begin
      CONVOLUTION_LOOP_for_for_for_x_lpi_1 <= MUX_v_8_2_2(z_out_5, CONVOLUTION_LOOP_for_for_for_for_asn_2929_mx0w0,
          CONVOLUTION_LOOP_for_for_for_for_for_and_5_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm <= {504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 504'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( core_wen & exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1_1 &
        main_stage_v_1 ) begin
      COMPUTE_LOOP_buf_tmp_lin_data_lpi_1_dfm <= buf_linear_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm <= {784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( core_wen & exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_1 & main_stage_v_1
        ) begin
      COMPUTE_LOOP_plm_tmp_f_data_lpi_1_dfm <= plm_kernel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_LOOP_asn_itm_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_74 | COMPUTE_LOOP_asn_itm_1_mx0c1) ) begin
      COMPUTE_LOOP_asn_itm_1 <= MUX_s_1_2_2(exit_COMPUTE_LOOP_lpi_1_dfm_3_mx0w0,
          exitL_exit_COMPUTE_LOOP_sva, COMPUTE_LOOP_asn_itm_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_74 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
          <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_25 & main_stage_v_1) | CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1)
        ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
          <= MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_sva_2_mx0w0, CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm,
          CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_3_st_1 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_42) ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_3_st_1 <= exit_COMPUTE_LOOP_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_8 & main_stage_v_2) | main_stage_v_3_mx0c1) )
        begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_3_st_2 <= 1'b0;
    end
    else if ( core_wen & (~(and_6_cse | and_dcpl_13 | (~ main_stage_v_2))) ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_3_st_2 <= exit_COMPUTE_LOOP_lpi_1_dfm_3_st_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_6_0_lpi_1_dfm <= 7'b0000000;
    end
    else if ( core_wen & main_stage_v_1 & exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1
        ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_6_0_lpi_1_dfm <= CONVOLUTION_LOOP_for_for_for_for_asn_2926_mx0w0;
    end
  end
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl = MUX_s_1_324_2(COMPUTE_LOOP_buf_tmp_acc_data_0_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_0_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_0_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_1_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_1_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_2_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_2_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_3_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_3_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_4_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_4_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_5_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_5_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_6_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_6_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_7_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_7_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_8_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_8_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_9_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_9_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_10_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_10_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_11_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_11_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_12_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_12_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_13_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_13_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_14_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_14_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_15_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_15_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_16_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_16_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_tmp_acc_data_17_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_tmp_acc_data_17_17_0_lpi_1_dfm_1_mx0, {CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1
      , (CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0]) , (CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1[0])});
  assign CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl = ~(MUX_v_30_2_2((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_tmp_acc_data_57_56_0_sat_sva_55_1_1[29:0]),
      30'b111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1));
  assign and_159_nl = exitL_exit_COMPUTE_LOOP_sva & and_tmp_14;
  assign or_135_nl = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)
      | (operator_8_false_1_acc_tmp[8]) | not_tmp_46;
  assign mux_46_nl = MUX_s_1_2_2(not_tmp_46, or_135_nl, operator_8_false_6_acc_itm_3_1);
  assign nand_26_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_42_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8])
      | not_tmp_46)));
  assign mux_47_nl = MUX_s_1_2_2(mux_46_nl, nand_26_nl, operator_8_false_5_acc_itm_3_1);
  assign and_149_nl = or_59_cse & or_155_cse & or_157_cse & nand_52_cse & nand_74_cse
      & (~((~(nor_32_cse | (CONVOLUTION_LOOP_for_acc_tmp[5]))) | mux_47_nl));
  assign mux_48_nl = MUX_s_1_2_2(and_159_nl, and_149_nl, main_stage_v_1);
  assign or_184_nl = CONVOLUTION_LOOP_for_for_if_CONVOLUTION_LOOP_for_for_if_nand_tmp
      | (operator_8_false_5_acc_tmp[8]) | nand_tmp_20;
  assign mux_62_nl = MUX_s_1_2_2(nand_tmp_20, or_184_nl, operator_8_false_3_acc_itm_4_1);
  assign mux_63_nl = MUX_s_1_2_2(and_tmp_29, (~ mux_62_nl), main_stage_v_1);
  assign mux_73_nl = MUX_s_1_2_2(and_tmp_29, (~ nand_tmp_20), main_stage_v_1);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_4_nl = MUX_v_3_2_2(CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2,
      ({{2{exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0}}, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0}),
      exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_1_dfm_1);
  assign CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_not_nl
      = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_for_not_26_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_not_339_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_1;
  assign CONVOLUTION_LOOP_for_for_not_14_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1;
  assign COMPUTE_LOOP_not_19_nl = ~ exitL_exit_COMPUTE_LOOP_sva_mx0;
  assign CONVOLUTION_LOOP_CONVOLUTION_LOOP_CONVOLUTION_LOOP_mux_nl = MUX_v_5_2_2((CONVOLUTION_LOOP_acc_tmp[4:0]),
      ({{4{or_155_cse}}, or_155_cse}), exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0);
  assign COMPUTE_LOOP_COMPUTE_LOOP_COMPUTE_LOOP_COMPUTE_LOOP_not_1_nl = ~ exitL_exit_COMPUTE_LOOP_sva_mx0;
  assign CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_mux_nl =
      MUX_v_5_2_2((CONVOLUTION_LOOP_for_acc_tmp[4:0]), ({{4{or_157_cse}}, or_157_cse}),
      exit_CONVOLUTION_LOOP_for_lpi_1_dfm_2_mx0);
  assign CONVOLUTION_LOOP_for_for_for_for_not_22_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
  assign operator_8_false_2_mux_4_nl = MUX_v_2_2_2((CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[1:0]),
      (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[4:3]), conf_info_crt_lpi_1_dfm_103_96_mx0[1]);
  assign operator_8_false_2_and_1_nl = (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[2])
      & (conf_info_crt_lpi_1_dfm_103_96_mx0[1]);
  assign operator_8_false_2_mux_5_nl = MUX_v_2_2_2((~ (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[3:2])),
      (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[7:6]), conf_info_crt_lpi_1_dfm_103_96_mx0[1]);
  assign nl_acc_nl = conv_u2u_3_4({operator_8_false_2_mux_4_nl , operator_8_false_2_and_1_nl})
      + conv_u2u_3_4({operator_8_false_2_mux_5_nl , 1'b1});
  assign acc_nl = nl_acc_nl[3:0];
  assign z_out = readslicef_4_3_1(acc_nl);
  assign operator_8_false_1_mux_2_nl = MUX_s_1_2_2((~ (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[1])),
      (~ (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[2])), conf_info_crt_lpi_1_dfm_103_96_mx0[2]);
  assign operator_8_false_1_and_1_nl = (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[6])
      & (~ (conf_info_crt_lpi_1_dfm_103_96_mx0[2]));
  assign operator_8_false_1_mux_3_nl = MUX_s_1_2_2((CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[2]),
      (~ (CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0[5])), conf_info_crt_lpi_1_dfm_103_96_mx0[2]);
  assign nl_acc_1_nl = conv_u2u_2_3({operator_8_false_1_mux_2_nl , operator_8_false_1_and_1_nl})
      + conv_u2u_2_3({operator_8_false_1_mux_3_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[2:0];
  assign z_out_1 = readslicef_3_2_1(acc_1_nl);
  assign nl_operator_8_false_3_acc_7_nl = ({(~ (operator_8_false_3_acc_imod_sva_1[2]))
      , 2'b00}) + conv_s2u_2_3(operator_8_false_3_acc_imod_sva_1[4:3]) + conv_u2u_1_3(operator_8_false_3_acc_imod_sva_1[2]);
  assign operator_8_false_3_acc_7_nl = nl_operator_8_false_3_acc_7_nl[2:0];
  assign operator_8_false_2_mux_6_nl = MUX_v_3_2_2(({(operator_8_false_2_acc_psp_1[2])
      , (operator_8_false_2_acc_psp_1[0]) , (operator_8_false_2_acc_5_sdt_1[0])}),
      operator_8_false_3_acc_7_nl, conf_info_crt_lpi_1_dfm_103_96_mx0[1]);
  assign nl_operator_8_false_2_acc_7_nl = conv_s2s_1_2(~ (operator_8_false_2_acc_psp_1[2]))
      + conv_u2s_1_2(~ (operator_8_false_2_acc_psp_1[1]));
  assign operator_8_false_2_acc_7_nl = nl_operator_8_false_2_acc_7_nl[1:0];
  assign operator_8_false_2_mux_7_nl = MUX_v_3_2_2((signext_3_2(operator_8_false_2_acc_7_nl)),
      ({1'b1 , (operator_8_false_3_acc_imod_sva_1[1:0])}), conf_info_crt_lpi_1_dfm_103_96_mx0[1]);
  assign nl_z_out_2_2_0 = operator_8_false_2_mux_6_nl + operator_8_false_2_mux_7_nl;
  assign z_out_2_2_0 = nl_z_out_2_2_0[2:0];
  assign nand_85_nl = ~((~((operator_8_false_1_acc_tmp[8:3]==6'b000000) & CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp))
      & operator_8_false_6_acc_itm_3_1);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_9_nl = MUX_v_8_2_2(({1'b0 , CONVOLUTION_LOOP_for_for_for_y_6_0_lpi_1_dfm_mx0}),
      CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0, nand_85_nl);
  assign nl_z_out_5 = CONVOLUTION_LOOP_for_for_for_for_for_mux_9_nl + 8'b00000001;
  assign z_out_5 = nl_z_out_5[7:0];

  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [54:0] MUX1HOT_v_55_3_2;
    input [54:0] input_2;
    input [54:0] input_1;
    input [54:0] input_0;
    input [2:0] sel;
    reg [54:0] result;
  begin
    result = input_0 & {55{sel[0]}};
    result = result | ( input_1 & {55{sel[1]}});
    result = result | ( input_2 & {55{sel[2]}});
    MUX1HOT_v_55_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_324_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] input_2;
    input [0:0] input_3;
    input [0:0] input_4;
    input [0:0] input_5;
    input [0:0] input_6;
    input [0:0] input_7;
    input [0:0] input_8;
    input [0:0] input_9;
    input [0:0] input_10;
    input [0:0] input_11;
    input [0:0] input_12;
    input [0:0] input_13;
    input [0:0] input_14;
    input [0:0] input_15;
    input [0:0] input_16;
    input [0:0] input_17;
    input [0:0] input_18;
    input [0:0] input_19;
    input [0:0] input_20;
    input [0:0] input_21;
    input [0:0] input_22;
    input [0:0] input_23;
    input [0:0] input_24;
    input [0:0] input_25;
    input [0:0] input_26;
    input [0:0] input_27;
    input [0:0] input_28;
    input [0:0] input_29;
    input [0:0] input_30;
    input [0:0] input_31;
    input [0:0] input_32;
    input [0:0] input_33;
    input [0:0] input_34;
    input [0:0] input_35;
    input [0:0] input_36;
    input [0:0] input_37;
    input [0:0] input_38;
    input [0:0] input_39;
    input [0:0] input_40;
    input [0:0] input_41;
    input [0:0] input_42;
    input [0:0] input_43;
    input [0:0] input_44;
    input [0:0] input_45;
    input [0:0] input_46;
    input [0:0] input_47;
    input [0:0] input_48;
    input [0:0] input_49;
    input [0:0] input_50;
    input [0:0] input_51;
    input [0:0] input_52;
    input [0:0] input_53;
    input [0:0] input_54;
    input [0:0] input_55;
    input [0:0] input_56;
    input [0:0] input_57;
    input [0:0] input_58;
    input [0:0] input_59;
    input [0:0] input_60;
    input [0:0] input_61;
    input [0:0] input_62;
    input [0:0] input_63;
    input [0:0] input_64;
    input [0:0] input_65;
    input [0:0] input_66;
    input [0:0] input_67;
    input [0:0] input_68;
    input [0:0] input_69;
    input [0:0] input_70;
    input [0:0] input_71;
    input [0:0] input_72;
    input [0:0] input_73;
    input [0:0] input_74;
    input [0:0] input_75;
    input [0:0] input_76;
    input [0:0] input_77;
    input [0:0] input_78;
    input [0:0] input_79;
    input [0:0] input_80;
    input [0:0] input_81;
    input [0:0] input_82;
    input [0:0] input_83;
    input [0:0] input_84;
    input [0:0] input_85;
    input [0:0] input_86;
    input [0:0] input_87;
    input [0:0] input_88;
    input [0:0] input_89;
    input [0:0] input_90;
    input [0:0] input_91;
    input [0:0] input_92;
    input [0:0] input_93;
    input [0:0] input_94;
    input [0:0] input_95;
    input [0:0] input_96;
    input [0:0] input_97;
    input [0:0] input_98;
    input [0:0] input_99;
    input [0:0] input_100;
    input [0:0] input_101;
    input [0:0] input_102;
    input [0:0] input_103;
    input [0:0] input_104;
    input [0:0] input_105;
    input [0:0] input_106;
    input [0:0] input_107;
    input [0:0] input_108;
    input [0:0] input_109;
    input [0:0] input_110;
    input [0:0] input_111;
    input [0:0] input_112;
    input [0:0] input_113;
    input [0:0] input_114;
    input [0:0] input_115;
    input [0:0] input_116;
    input [0:0] input_117;
    input [0:0] input_118;
    input [0:0] input_119;
    input [0:0] input_120;
    input [0:0] input_121;
    input [0:0] input_122;
    input [0:0] input_123;
    input [0:0] input_124;
    input [0:0] input_125;
    input [0:0] input_126;
    input [0:0] input_127;
    input [0:0] input_128;
    input [0:0] input_129;
    input [0:0] input_130;
    input [0:0] input_131;
    input [0:0] input_132;
    input [0:0] input_133;
    input [0:0] input_134;
    input [0:0] input_135;
    input [0:0] input_136;
    input [0:0] input_137;
    input [0:0] input_138;
    input [0:0] input_139;
    input [0:0] input_140;
    input [0:0] input_141;
    input [0:0] input_142;
    input [0:0] input_143;
    input [0:0] input_144;
    input [0:0] input_145;
    input [0:0] input_146;
    input [0:0] input_147;
    input [0:0] input_148;
    input [0:0] input_149;
    input [0:0] input_150;
    input [0:0] input_151;
    input [0:0] input_152;
    input [0:0] input_153;
    input [0:0] input_154;
    input [0:0] input_155;
    input [0:0] input_156;
    input [0:0] input_157;
    input [0:0] input_158;
    input [0:0] input_159;
    input [0:0] input_160;
    input [0:0] input_161;
    input [0:0] input_162;
    input [0:0] input_163;
    input [0:0] input_164;
    input [0:0] input_165;
    input [0:0] input_166;
    input [0:0] input_167;
    input [0:0] input_168;
    input [0:0] input_169;
    input [0:0] input_170;
    input [0:0] input_171;
    input [0:0] input_172;
    input [0:0] input_173;
    input [0:0] input_174;
    input [0:0] input_175;
    input [0:0] input_176;
    input [0:0] input_177;
    input [0:0] input_178;
    input [0:0] input_179;
    input [0:0] input_180;
    input [0:0] input_181;
    input [0:0] input_182;
    input [0:0] input_183;
    input [0:0] input_184;
    input [0:0] input_185;
    input [0:0] input_186;
    input [0:0] input_187;
    input [0:0] input_188;
    input [0:0] input_189;
    input [0:0] input_190;
    input [0:0] input_191;
    input [0:0] input_192;
    input [0:0] input_193;
    input [0:0] input_194;
    input [0:0] input_195;
    input [0:0] input_196;
    input [0:0] input_197;
    input [0:0] input_198;
    input [0:0] input_199;
    input [0:0] input_200;
    input [0:0] input_201;
    input [0:0] input_202;
    input [0:0] input_203;
    input [0:0] input_204;
    input [0:0] input_205;
    input [0:0] input_206;
    input [0:0] input_207;
    input [0:0] input_208;
    input [0:0] input_209;
    input [0:0] input_210;
    input [0:0] input_211;
    input [0:0] input_212;
    input [0:0] input_213;
    input [0:0] input_214;
    input [0:0] input_215;
    input [0:0] input_216;
    input [0:0] input_217;
    input [0:0] input_218;
    input [0:0] input_219;
    input [0:0] input_220;
    input [0:0] input_221;
    input [0:0] input_222;
    input [0:0] input_223;
    input [0:0] input_224;
    input [0:0] input_225;
    input [0:0] input_226;
    input [0:0] input_227;
    input [0:0] input_228;
    input [0:0] input_229;
    input [0:0] input_230;
    input [0:0] input_231;
    input [0:0] input_232;
    input [0:0] input_233;
    input [0:0] input_234;
    input [0:0] input_235;
    input [0:0] input_236;
    input [0:0] input_237;
    input [0:0] input_238;
    input [0:0] input_239;
    input [0:0] input_240;
    input [0:0] input_241;
    input [0:0] input_242;
    input [0:0] input_243;
    input [0:0] input_244;
    input [0:0] input_245;
    input [0:0] input_246;
    input [0:0] input_247;
    input [0:0] input_248;
    input [0:0] input_249;
    input [0:0] input_250;
    input [0:0] input_251;
    input [0:0] input_252;
    input [0:0] input_253;
    input [0:0] input_254;
    input [0:0] input_255;
    input [0:0] input_256;
    input [0:0] input_257;
    input [0:0] input_258;
    input [0:0] input_259;
    input [0:0] input_260;
    input [0:0] input_261;
    input [0:0] input_262;
    input [0:0] input_263;
    input [0:0] input_264;
    input [0:0] input_265;
    input [0:0] input_266;
    input [0:0] input_267;
    input [0:0] input_268;
    input [0:0] input_269;
    input [0:0] input_270;
    input [0:0] input_271;
    input [0:0] input_272;
    input [0:0] input_273;
    input [0:0] input_274;
    input [0:0] input_275;
    input [0:0] input_276;
    input [0:0] input_277;
    input [0:0] input_278;
    input [0:0] input_279;
    input [0:0] input_280;
    input [0:0] input_281;
    input [0:0] input_282;
    input [0:0] input_283;
    input [0:0] input_284;
    input [0:0] input_285;
    input [0:0] input_286;
    input [0:0] input_287;
    input [0:0] input_288;
    input [0:0] input_289;
    input [0:0] input_290;
    input [0:0] input_291;
    input [0:0] input_292;
    input [0:0] input_293;
    input [0:0] input_294;
    input [0:0] input_295;
    input [0:0] input_296;
    input [0:0] input_297;
    input [0:0] input_298;
    input [0:0] input_299;
    input [0:0] input_300;
    input [0:0] input_301;
    input [0:0] input_302;
    input [0:0] input_303;
    input [0:0] input_304;
    input [0:0] input_305;
    input [0:0] input_306;
    input [0:0] input_307;
    input [0:0] input_308;
    input [0:0] input_309;
    input [0:0] input_310;
    input [0:0] input_311;
    input [0:0] input_312;
    input [0:0] input_313;
    input [0:0] input_314;
    input [0:0] input_315;
    input [0:0] input_316;
    input [0:0] input_317;
    input [0:0] input_318;
    input [0:0] input_319;
    input [0:0] input_320;
    input [0:0] input_321;
    input [0:0] input_322;
    input [0:0] input_323;
    input [8:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_s_1_324_2 = result;
  end
  endfunction


  function automatic [1567:0] MUX_v_1568_2_2;
    input [1567:0] input_0;
    input [1567:0] input_1;
    input [0:0] sel;
    reg [1567:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_1568_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_126_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [31:0] input_32;
    input [31:0] input_33;
    input [31:0] input_34;
    input [31:0] input_35;
    input [31:0] input_36;
    input [31:0] input_37;
    input [31:0] input_38;
    input [31:0] input_39;
    input [31:0] input_40;
    input [31:0] input_41;
    input [31:0] input_42;
    input [31:0] input_43;
    input [31:0] input_44;
    input [31:0] input_45;
    input [31:0] input_46;
    input [31:0] input_47;
    input [31:0] input_48;
    input [31:0] input_49;
    input [31:0] input_50;
    input [31:0] input_51;
    input [31:0] input_52;
    input [31:0] input_53;
    input [31:0] input_54;
    input [31:0] input_55;
    input [31:0] input_56;
    input [31:0] input_57;
    input [31:0] input_58;
    input [31:0] input_59;
    input [31:0] input_60;
    input [31:0] input_61;
    input [31:0] input_62;
    input [31:0] input_63;
    input [31:0] input_64;
    input [31:0] input_65;
    input [31:0] input_66;
    input [31:0] input_67;
    input [31:0] input_68;
    input [31:0] input_69;
    input [31:0] input_70;
    input [31:0] input_71;
    input [31:0] input_72;
    input [31:0] input_73;
    input [31:0] input_74;
    input [31:0] input_75;
    input [31:0] input_76;
    input [31:0] input_77;
    input [31:0] input_78;
    input [31:0] input_79;
    input [31:0] input_80;
    input [31:0] input_81;
    input [31:0] input_82;
    input [31:0] input_83;
    input [31:0] input_84;
    input [31:0] input_85;
    input [31:0] input_86;
    input [31:0] input_87;
    input [31:0] input_88;
    input [31:0] input_89;
    input [31:0] input_90;
    input [31:0] input_91;
    input [31:0] input_92;
    input [31:0] input_93;
    input [31:0] input_94;
    input [31:0] input_95;
    input [31:0] input_96;
    input [31:0] input_97;
    input [31:0] input_98;
    input [31:0] input_99;
    input [31:0] input_100;
    input [31:0] input_101;
    input [31:0] input_102;
    input [31:0] input_103;
    input [31:0] input_104;
    input [31:0] input_105;
    input [31:0] input_106;
    input [31:0] input_107;
    input [31:0] input_108;
    input [31:0] input_109;
    input [31:0] input_110;
    input [31:0] input_111;
    input [31:0] input_112;
    input [31:0] input_113;
    input [31:0] input_114;
    input [31:0] input_115;
    input [31:0] input_116;
    input [31:0] input_117;
    input [31:0] input_118;
    input [31:0] input_119;
    input [31:0] input_120;
    input [31:0] input_121;
    input [31:0] input_122;
    input [31:0] input_123;
    input [31:0] input_124;
    input [31:0] input_125;
    input [6:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      default : begin
        result = input_125;
      end
    endcase
    MUX_v_32_126_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_49_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [31:0] input_32;
    input [31:0] input_33;
    input [31:0] input_34;
    input [31:0] input_35;
    input [31:0] input_36;
    input [31:0] input_37;
    input [31:0] input_38;
    input [31:0] input_39;
    input [31:0] input_40;
    input [31:0] input_41;
    input [31:0] input_42;
    input [31:0] input_43;
    input [31:0] input_44;
    input [31:0] input_45;
    input [31:0] input_46;
    input [31:0] input_47;
    input [31:0] input_48;
    input [5:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      default : begin
        result = input_48;
      end
    endcase
    MUX_v_32_49_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [4031:0] MUX_v_4032_2_2;
    input [4031:0] input_0;
    input [4031:0] input_1;
    input [0:0] sel;
    reg [4031:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4032_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [54:0] MUX_v_55_2_2;
    input [54:0] input_0;
    input [54:0] input_1;
    input [0:0] sel;
    reg [54:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_55_2_2 = result;
  end
  endfunction


  function automatic [54:0] MUX_v_55_324_2;
    input [54:0] input_0;
    input [54:0] input_1;
    input [54:0] input_2;
    input [54:0] input_3;
    input [54:0] input_4;
    input [54:0] input_5;
    input [54:0] input_6;
    input [54:0] input_7;
    input [54:0] input_8;
    input [54:0] input_9;
    input [54:0] input_10;
    input [54:0] input_11;
    input [54:0] input_12;
    input [54:0] input_13;
    input [54:0] input_14;
    input [54:0] input_15;
    input [54:0] input_16;
    input [54:0] input_17;
    input [54:0] input_18;
    input [54:0] input_19;
    input [54:0] input_20;
    input [54:0] input_21;
    input [54:0] input_22;
    input [54:0] input_23;
    input [54:0] input_24;
    input [54:0] input_25;
    input [54:0] input_26;
    input [54:0] input_27;
    input [54:0] input_28;
    input [54:0] input_29;
    input [54:0] input_30;
    input [54:0] input_31;
    input [54:0] input_32;
    input [54:0] input_33;
    input [54:0] input_34;
    input [54:0] input_35;
    input [54:0] input_36;
    input [54:0] input_37;
    input [54:0] input_38;
    input [54:0] input_39;
    input [54:0] input_40;
    input [54:0] input_41;
    input [54:0] input_42;
    input [54:0] input_43;
    input [54:0] input_44;
    input [54:0] input_45;
    input [54:0] input_46;
    input [54:0] input_47;
    input [54:0] input_48;
    input [54:0] input_49;
    input [54:0] input_50;
    input [54:0] input_51;
    input [54:0] input_52;
    input [54:0] input_53;
    input [54:0] input_54;
    input [54:0] input_55;
    input [54:0] input_56;
    input [54:0] input_57;
    input [54:0] input_58;
    input [54:0] input_59;
    input [54:0] input_60;
    input [54:0] input_61;
    input [54:0] input_62;
    input [54:0] input_63;
    input [54:0] input_64;
    input [54:0] input_65;
    input [54:0] input_66;
    input [54:0] input_67;
    input [54:0] input_68;
    input [54:0] input_69;
    input [54:0] input_70;
    input [54:0] input_71;
    input [54:0] input_72;
    input [54:0] input_73;
    input [54:0] input_74;
    input [54:0] input_75;
    input [54:0] input_76;
    input [54:0] input_77;
    input [54:0] input_78;
    input [54:0] input_79;
    input [54:0] input_80;
    input [54:0] input_81;
    input [54:0] input_82;
    input [54:0] input_83;
    input [54:0] input_84;
    input [54:0] input_85;
    input [54:0] input_86;
    input [54:0] input_87;
    input [54:0] input_88;
    input [54:0] input_89;
    input [54:0] input_90;
    input [54:0] input_91;
    input [54:0] input_92;
    input [54:0] input_93;
    input [54:0] input_94;
    input [54:0] input_95;
    input [54:0] input_96;
    input [54:0] input_97;
    input [54:0] input_98;
    input [54:0] input_99;
    input [54:0] input_100;
    input [54:0] input_101;
    input [54:0] input_102;
    input [54:0] input_103;
    input [54:0] input_104;
    input [54:0] input_105;
    input [54:0] input_106;
    input [54:0] input_107;
    input [54:0] input_108;
    input [54:0] input_109;
    input [54:0] input_110;
    input [54:0] input_111;
    input [54:0] input_112;
    input [54:0] input_113;
    input [54:0] input_114;
    input [54:0] input_115;
    input [54:0] input_116;
    input [54:0] input_117;
    input [54:0] input_118;
    input [54:0] input_119;
    input [54:0] input_120;
    input [54:0] input_121;
    input [54:0] input_122;
    input [54:0] input_123;
    input [54:0] input_124;
    input [54:0] input_125;
    input [54:0] input_126;
    input [54:0] input_127;
    input [54:0] input_128;
    input [54:0] input_129;
    input [54:0] input_130;
    input [54:0] input_131;
    input [54:0] input_132;
    input [54:0] input_133;
    input [54:0] input_134;
    input [54:0] input_135;
    input [54:0] input_136;
    input [54:0] input_137;
    input [54:0] input_138;
    input [54:0] input_139;
    input [54:0] input_140;
    input [54:0] input_141;
    input [54:0] input_142;
    input [54:0] input_143;
    input [54:0] input_144;
    input [54:0] input_145;
    input [54:0] input_146;
    input [54:0] input_147;
    input [54:0] input_148;
    input [54:0] input_149;
    input [54:0] input_150;
    input [54:0] input_151;
    input [54:0] input_152;
    input [54:0] input_153;
    input [54:0] input_154;
    input [54:0] input_155;
    input [54:0] input_156;
    input [54:0] input_157;
    input [54:0] input_158;
    input [54:0] input_159;
    input [54:0] input_160;
    input [54:0] input_161;
    input [54:0] input_162;
    input [54:0] input_163;
    input [54:0] input_164;
    input [54:0] input_165;
    input [54:0] input_166;
    input [54:0] input_167;
    input [54:0] input_168;
    input [54:0] input_169;
    input [54:0] input_170;
    input [54:0] input_171;
    input [54:0] input_172;
    input [54:0] input_173;
    input [54:0] input_174;
    input [54:0] input_175;
    input [54:0] input_176;
    input [54:0] input_177;
    input [54:0] input_178;
    input [54:0] input_179;
    input [54:0] input_180;
    input [54:0] input_181;
    input [54:0] input_182;
    input [54:0] input_183;
    input [54:0] input_184;
    input [54:0] input_185;
    input [54:0] input_186;
    input [54:0] input_187;
    input [54:0] input_188;
    input [54:0] input_189;
    input [54:0] input_190;
    input [54:0] input_191;
    input [54:0] input_192;
    input [54:0] input_193;
    input [54:0] input_194;
    input [54:0] input_195;
    input [54:0] input_196;
    input [54:0] input_197;
    input [54:0] input_198;
    input [54:0] input_199;
    input [54:0] input_200;
    input [54:0] input_201;
    input [54:0] input_202;
    input [54:0] input_203;
    input [54:0] input_204;
    input [54:0] input_205;
    input [54:0] input_206;
    input [54:0] input_207;
    input [54:0] input_208;
    input [54:0] input_209;
    input [54:0] input_210;
    input [54:0] input_211;
    input [54:0] input_212;
    input [54:0] input_213;
    input [54:0] input_214;
    input [54:0] input_215;
    input [54:0] input_216;
    input [54:0] input_217;
    input [54:0] input_218;
    input [54:0] input_219;
    input [54:0] input_220;
    input [54:0] input_221;
    input [54:0] input_222;
    input [54:0] input_223;
    input [54:0] input_224;
    input [54:0] input_225;
    input [54:0] input_226;
    input [54:0] input_227;
    input [54:0] input_228;
    input [54:0] input_229;
    input [54:0] input_230;
    input [54:0] input_231;
    input [54:0] input_232;
    input [54:0] input_233;
    input [54:0] input_234;
    input [54:0] input_235;
    input [54:0] input_236;
    input [54:0] input_237;
    input [54:0] input_238;
    input [54:0] input_239;
    input [54:0] input_240;
    input [54:0] input_241;
    input [54:0] input_242;
    input [54:0] input_243;
    input [54:0] input_244;
    input [54:0] input_245;
    input [54:0] input_246;
    input [54:0] input_247;
    input [54:0] input_248;
    input [54:0] input_249;
    input [54:0] input_250;
    input [54:0] input_251;
    input [54:0] input_252;
    input [54:0] input_253;
    input [54:0] input_254;
    input [54:0] input_255;
    input [54:0] input_256;
    input [54:0] input_257;
    input [54:0] input_258;
    input [54:0] input_259;
    input [54:0] input_260;
    input [54:0] input_261;
    input [54:0] input_262;
    input [54:0] input_263;
    input [54:0] input_264;
    input [54:0] input_265;
    input [54:0] input_266;
    input [54:0] input_267;
    input [54:0] input_268;
    input [54:0] input_269;
    input [54:0] input_270;
    input [54:0] input_271;
    input [54:0] input_272;
    input [54:0] input_273;
    input [54:0] input_274;
    input [54:0] input_275;
    input [54:0] input_276;
    input [54:0] input_277;
    input [54:0] input_278;
    input [54:0] input_279;
    input [54:0] input_280;
    input [54:0] input_281;
    input [54:0] input_282;
    input [54:0] input_283;
    input [54:0] input_284;
    input [54:0] input_285;
    input [54:0] input_286;
    input [54:0] input_287;
    input [54:0] input_288;
    input [54:0] input_289;
    input [54:0] input_290;
    input [54:0] input_291;
    input [54:0] input_292;
    input [54:0] input_293;
    input [54:0] input_294;
    input [54:0] input_295;
    input [54:0] input_296;
    input [54:0] input_297;
    input [54:0] input_298;
    input [54:0] input_299;
    input [54:0] input_300;
    input [54:0] input_301;
    input [54:0] input_302;
    input [54:0] input_303;
    input [54:0] input_304;
    input [54:0] input_305;
    input [54:0] input_306;
    input [54:0] input_307;
    input [54:0] input_308;
    input [54:0] input_309;
    input [54:0] input_310;
    input [54:0] input_311;
    input [54:0] input_312;
    input [54:0] input_313;
    input [54:0] input_314;
    input [54:0] input_315;
    input [54:0] input_316;
    input [54:0] input_317;
    input [54:0] input_318;
    input [54:0] input_319;
    input [54:0] input_320;
    input [54:0] input_321;
    input [54:0] input_322;
    input [54:0] input_323;
    input [8:0] sel;
    reg [54:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_v_55_324_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [1:0] readslicef_3_2_1;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_3_2_1 = tmp[1:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [2:0] readslicef_4_3_1;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_4_3_1 = tmp[2:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function automatic [2:0] signext_3_2;
    input [1:0] vector;
  begin
    signext_3_2= {{1{vector[1]}}, vector};
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [2:0] conv_s2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_3 = {vector[1], vector};
  end
  endfunction


  function automatic [3:0] conv_s2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2s_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_9_17 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_17 = {{8{vector[8]}}, vector};
  end
  endfunction


  function automatic [57:0] conv_s2s_57_58 ;
    input [56:0]  vector ;
  begin
    conv_s2s_57_58 = {vector[56], vector};
  end
  endfunction


  function automatic [2:0] conv_s2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_3 = {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] conv_s2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_3 = {vector[1], vector};
  end
  endfunction


  function automatic [57:0] conv_s2u_48_58 ;
    input [47:0]  vector ;
  begin
    conv_s2u_48_58 = {{10{vector[47]}}, vector};
  end
  endfunction


  function automatic [57:0] conv_s2u_57_58 ;
    input [56:0]  vector ;
  begin
    conv_s2u_57_58 = {vector[56], vector};
  end
  endfunction


  function automatic [63:0] conv_s2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_s2u_64_64 = vector;
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [57:0] conv_u2s_1_58 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_58 = {{57{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_3 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_2_5 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_5 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_3_6 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_6 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store_core
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, var_output_rsc_dat,
      var_output_rsc_vld, var_output_rsc_rdy, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld,
      dma_write_ctrl_rsc_rdy, dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input [31:0] var_output_rsc_dat;
  input var_output_rsc_vld;
  output var_output_rsc_rdy;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire core_wen;
  wire conf_info_rsci_bawt;
  wire conf_info_rsci_wen_comp;
  wire [63:0] conf_info_rsci_idat_mxwt;
  wire var_output_rsci_bawt;
  wire var_output_rsci_wen_comp;
  wire [31:0] var_output_rsci_idat_mxwt;
  wire dma_write_ctrl_rsci_bawt;
  wire dma_write_ctrl_rsci_wen_comp;
  wire dma_write_chnl_rsci_bawt;
  wire dma_write_chnl_rsci_wen_comp;
  wire done_rsci_bawt;
  wire done_rsci_wen_comp;
  reg [15:0] dma_write_ctrl_rsci_idat_15_0;
  reg [31:0] dma_write_chnl_rsci_idat_31_0;
  wire [1:0] fsm_output;
  wire [8:0] operator_8_false_4_acc_tmp;
  wire [9:0] nl_operator_8_false_4_acc_tmp;
  wire [5:0] STORE_INNER_LOOP_acc_tmp;
  wire [6:0] nl_STORE_INNER_LOOP_acc_tmp;
  wire [8:0] operator_8_false_3_acc_tmp;
  wire [9:0] nl_operator_8_false_3_acc_tmp;
  wire [8:0] operator_8_false_2_acc_tmp;
  wire [9:0] nl_operator_8_false_2_acc_tmp;
  wire STORE_INNER_LOOP_for_for_if_1_STORE_INNER_LOOP_for_for_if_1_nand_tmp;
  wire [8:0] operator_8_false_1_acc_tmp;
  wire [9:0] nl_operator_8_false_1_acc_tmp;
  wire or_tmp_7;
  wire and_tmp_4;
  wire mux_tmp_16;
  wire and_tmp_5;
  wire mux_tmp_17;
  wire nand_tmp_4;
  wire or_tmp_40;
  wire nand_tmp_5;
  wire and_dcpl_9;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_30;
  wire and_dcpl_34;
  wire and_dcpl_42;
  wire and_dcpl_45;
  wire or_dcpl_20;
  wire or_dcpl_21;
  wire or_dcpl_22;
  wire or_dcpl_25;
  wire and_dcpl_46;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_56;
  wire or_dcpl_33;
  wire or_tmp_56;
  wire or_tmp_70;
  wire main_stage_en_3;
  wire [4:0] STORE_BATCH_LOOP_b_4_0_sva_2;
  wire [5:0] nl_STORE_BATCH_LOOP_b_4_0_sva_2;
  wire exit_STORE_INNER_LOOP_lpi_1_dfm_3_mx0w0;
  wire [3:0] STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1;
  wire exit_STORE_INNER_LOOP_for_lpi_1_dfm_3_mx0w0;
  wire [4:0] STORE_INNER_LOOP_fl_5_0_lpi_1_dfm_4_0_1;
  wire [4:0] STORE_INNER_LOOP_for_i_4_0_lpi_1_dfm_4;
  wire [4:0] STORE_INNER_LOOP_for_for_j_4_0_lpi_1_dfm_3;
  reg exit_STORE_INNER_LOOP_lpi_1_dfm_3;
  wire unequal_tmp_1;
  reg exitL_exit_STORE_BATCH_LOOP_sva;
  reg STORE_BATCH_LOOP_asn_itm;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2;
  reg main_stage_v_2;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1;
  wire exit_STORE_BATCH_LOOP_sva_2_mx0w0;
  reg exit_STORE_BATCH_LOOP_sva_2;
  reg exit_STORE_INNER_LOOP_lpi_1_dfm_1;
  wire exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0;
  reg exit_STORE_INNER_LOOP_for_lpi_1_dfm_1;
  reg reg_conf_info_rsci_iswt0_cse;
  wire STORE_BATCH_LOOP_and_2_cse;
  reg reg_done_rsci_ivld_core_psct_cse;
  reg reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  wire or_138_cse;
  wire nor_23_cse;
  wire or_64_cse;
  wire or_5_cse;
  wire and_165_cse;
  wire and_7_cse;
  wire or_139_cse;
  wire and_158_cse;
  wire or_59_cse;
  wire and_162_cse;
  wire or_57_cse;
  wire and_160_cse;
  wire [10:0] z_out;
  wire [10:0] z_out_1;
  wire [9:0] z_out_2;
  reg [15:0] dma_write_data_index_lpi_1;
  wire [16:0] nl_dma_write_data_index_lpi_1;
  reg [4:0] STORE_INNER_LOOP_for_i_4_0_lpi_1;
  reg [4:0] STORE_INNER_LOOP_for_for_j_4_0_lpi_1;
  reg [7:0] n_w_out_lpi_1_dfm_1;
  reg [7:0] n_h_out_lpi_1_dfm_1;
  reg exit_STORE_INNER_LOOP_for_lpi_1_dfm_3;
  reg [3:0] STORE_BATCH_LOOP_b_4_0_lpi_1_3_0;
  reg [4:0] STORE_INNER_LOOP_fl_5_0_lpi_1_4_0;
  reg [7:0] conf_info_crt_lpi_1_dfm_231_224;
  reg [7:0] conf_info_crt_lpi_1_dfm_199_192;
  reg [7:0] conf_info_crt_lpi_1_dfm_167_160;
  reg [7:0] conf_info_crt_lpi_1_dfm_135_128;
  reg [7:0] conf_info_crt_lpi_1_dfm_103_96;
  reg [7:0] conf_info_crt_lpi_1_dfm_71_64;
  wire [15:0] dma_write_data_index_lpi_1_dfm_mx1w0;
  wire [16:0] nl_dma_write_data_index_lpi_1_dfm_mx1w0;
  wire [7:0] conf_info_crt_lpi_1_dfm_199_192_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_167_160_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_135_128_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_103_96_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_71_64_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_231_224_mx0;
  wire [7:0] n_w_out_lpi_1_dfm_3;
  wire [7:0] n_h_out_lpi_1_dfm_3;
  wire exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
  wire main_stage_v_2_mx0c1;
  wire [7:0] pad_sva_1;
  wire signed [16:0] nl_pad_sva_1;
  wire [16:0] pad_acc_psp_sva_1;
  wire [17:0] nl_pad_acc_psp_sva_1;
  wire [4:0] STORE_INNER_LOOP_for_i_4_0_sva_2;
  wire [5:0] nl_STORE_INNER_LOOP_for_i_4_0_sva_2;
  wire [4:0] STORE_INNER_LOOP_for_for_j_4_0_sva_2;
  wire [5:0] nl_STORE_INNER_LOOP_for_for_j_4_0_sva_2;
  wire STORE_BATCH_LOOP_asn_41;
  wire STORE_BATCH_LOOP_asn_43;
  wire and_34_rgt;
  wire and_64_rgt;
  wire STORE_INNER_LOOP_for_and_3_rgt;
  wire STORE_INNER_LOOP_for_and_4_rgt;
  wire and_76_rgt;
  reg reg_var_output_rsci_iswt0_cse;
  wire and_185_cse;
  wire n_w_out_and_cse;
  wire mux_43_itm;
  wire operator_8_false_2_acc_itm_4_1;
  wire operator_8_false_3_acc_itm_4_1;
  wire [1:0] if_if_and_cse;
  wire if_if_nand_2_cse;

  wire[0:0] mux_26_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] mux_22_nl;
  wire[15:0] dma_write_data_index_mux_1_nl;
  wire[0:0] nor_41_nl;
  wire[0:0] and_18_nl;
  wire[0:0] mux_28_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_nl;
  wire[15:0] STORE_BATCH_LOOP_acc_1_nl;
  wire[16:0] nl_STORE_BATCH_LOOP_acc_1_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_1_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_1_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_2_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_3_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_3_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_4_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_4_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_5_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_6_nl;
  wire[19:0] nl_STORE_BATCH_LOOP_mul_6_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_7_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_7_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_8_nl;
  wire[7:0] operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_acc_nl;
  wire[0:0] operator_42_true_and_nl;
  wire[7:0] operator_43_true_1_acc_nl;
  wire[8:0] nl_operator_43_true_1_acc_nl;
  wire[0:0] operator_42_true_1_and_nl;
  wire[0:0] STORE_BATCH_LOOP_mux_8_nl;
  wire[0:0] or_83_nl;
  wire[0:0] STORE_INNER_LOOP_mux_1_nl;
  wire[0:0] STORE_INNER_LOOP_for_mux_1_nl;
  wire[7:0] operator_43_true_operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_operator_43_true_acc_nl;
  wire[0:0] operator_43_true_and_nl;
  wire[8:0] pad_acc_2_nl;
  wire[9:0] nl_pad_acc_2_nl;
  wire[16:0] pad_mul_nl;
  wire signed [17:0] nl_pad_mul_nl;
  wire[8:0] operator_8_false_acc_nl;
  wire[9:0] nl_operator_8_false_acc_nl;
  wire[0:0] STORE_BATCH_LOOP_not_27_nl;
  wire[0:0] STORE_INNER_LOOP_not_14_nl;
  wire[4:0] operator_8_false_2_acc_nl;
  wire[5:0] nl_operator_8_false_2_acc_nl;
  wire[0:0] STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_BATCH_LOOP_not_nl;
  wire[4:0] operator_8_false_3_acc_nl;
  wire[5:0] nl_operator_8_false_3_acc_nl;
  wire[0:0] STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_INNER_LOOP_nor_nl;
  wire[0:0] nor_42_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] or_89_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] mux_44_nl;
  wire[11:0] acc_nl;
  wire[12:0] nl_acc_nl;
  wire[11:0] acc_1_nl;
  wire[12:0] nl_acc_1_nl;
  wire[10:0] acc_2_nl;
  wire[11:0] nl_acc_2_nl;
  wire[0:0] if_if_and_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_store_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg;
  assign nl_store_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg = conf_info_rsci_bawt
      & STORE_BATCH_LOOP_asn_itm & var_output_rsci_bawt & mux_tmp_16 & (fsm_output[1]);
  wire [66:0] nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat;
  assign nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat = {51'b011000000000000000000000000000000010000000000000000
      , dma_write_ctrl_rsci_idat_15_0};
  wire [63:0] nl_store_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat;
  assign nl_store_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat = {32'b11011110101011011011111011101111
      , dma_write_chnl_rsci_idat_31_0};
  esp_acc_conv2dlb_cxx_catapult_store_core_conf_info_rsci store_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(nl_store_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg[0:0]),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_iswt0(reg_conf_info_rsci_iswt0_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_var_output_rsci store_core_var_output_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .var_output_rsc_dat(var_output_rsc_dat),
      .var_output_rsc_vld(var_output_rsc_vld),
      .var_output_rsc_rdy(var_output_rsc_rdy),
      .core_wen(core_wen),
      .var_output_rsci_oswt_unreg(or_tmp_70),
      .var_output_rsci_bawt(var_output_rsci_bawt),
      .var_output_rsci_iswt0(reg_var_output_rsci_iswt0_cse),
      .var_output_rsci_wen_comp(var_output_rsci_wen_comp),
      .var_output_rsci_idat_mxwt(var_output_rsci_idat_mxwt)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_ctrl_rsci store_core_dma_write_ctrl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .core_wen(core_wen),
      .dma_write_ctrl_rsci_oswt_unreg(and_dcpl_34),
      .dma_write_ctrl_rsci_bawt(dma_write_ctrl_rsci_bawt),
      .dma_write_ctrl_rsci_iswt0(reg_dma_write_chnl_rsci_ivld_core_psct_cse),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_ctrl_rsci_idat(nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat[66:0])
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_dma_write_chnl_rsci store_core_dma_write_chnl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .core_wen(core_wen),
      .dma_write_chnl_rsci_oswt_unreg(and_dcpl_34),
      .dma_write_chnl_rsci_bawt(dma_write_chnl_rsci_bawt),
      .dma_write_chnl_rsci_iswt0(reg_dma_write_chnl_rsci_ivld_core_psct_cse),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .dma_write_chnl_rsci_idat(nl_store_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat[63:0])
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_done_rsci store_core_done_rsci_inst (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(and_dcpl_26),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_iswt0(reg_done_rsci_ivld_core_psct_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_staller store_core_staller_inst (
      .core_wen(core_wen),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .var_output_rsci_wen_comp(var_output_rsci_wen_comp),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2dlb_cxx_catapult_store_core_core_fsm store_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_158_cse = or_139_cse & operator_8_false_2_acc_itm_4_1;
  assign or_59_cse = nor_23_cse | (STORE_INNER_LOOP_acc_tmp[5]);
  assign or_57_cse = exit_STORE_BATCH_LOOP_sva_2_mx0w0 | (STORE_BATCH_LOOP_b_4_0_sva_2[4]);
  assign STORE_BATCH_LOOP_and_2_cse = core_wen & (~((~ mux_tmp_17) | (fsm_output[0])));
  assign or_64_cse = exitL_exit_STORE_BATCH_LOOP_sva | exit_STORE_INNER_LOOP_lpi_1_dfm_3
      | exit_STORE_BATCH_LOOP_lpi_1_dfm_2;
  assign or_5_cse = (~ STORE_BATCH_LOOP_asn_itm) | conf_info_rsci_bawt;
  assign and_34_rgt = and_dcpl_9 & var_output_rsci_bawt & (~ exitL_exit_STORE_BATCH_LOOP_sva)
      & (~ exit_STORE_INNER_LOOP_lpi_1_dfm_3) & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_2);
  assign and_160_cse = or_5_cse & var_output_rsci_bawt;
  assign n_w_out_and_cse = core_wen & mux_tmp_17;
  assign or_138_cse = STORE_INNER_LOOP_for_for_if_1_STORE_INNER_LOOP_for_for_if_1_nand_tmp
      | (operator_8_false_1_acc_tmp[8]);
  assign or_139_cse = (~((STORE_INNER_LOOP_for_i_4_0_lpi_1_dfm_4 == (operator_8_false_2_acc_tmp[4:0]))
      & (operator_8_false_2_acc_tmp[7:5]==3'b000))) | (operator_8_false_2_acc_tmp[8]);
  assign and_162_cse = or_138_cse & operator_8_false_3_acc_itm_4_1;
  assign and_64_rgt = and_dcpl_9 & or_138_cse & var_output_rsci_bawt & operator_8_false_3_acc_itm_4_1;
  assign STORE_INNER_LOOP_for_and_3_rgt = (~ and_162_cse) & and_dcpl_56;
  assign STORE_INNER_LOOP_for_and_4_rgt = and_162_cse & and_dcpl_56;
  assign nor_23_cse = ~((operator_8_false_3_acc_tmp[8]) | (~((STORE_INNER_LOOP_fl_5_0_lpi_1_dfm_4_0_1
      == (operator_8_false_3_acc_tmp[4:0])) & (operator_8_false_3_acc_tmp[7:5]==3'b000))));
  assign and_18_nl = operator_8_false_3_acc_itm_4_1 & or_138_cse & nand_tmp_5;
  assign mux_43_itm = MUX_s_1_2_2(and_18_nl, nand_tmp_5, and_158_cse);
  assign mux_28_nl = MUX_s_1_2_2(nand_tmp_5, mux_43_itm, or_59_cse);
  assign and_76_rgt = mux_28_nl & or_tmp_7 & and_160_cse;
  assign STORE_BATCH_LOOP_mul_2_nl = conv_u2u_16_16(conf_info_crt_lpi_1_dfm_199_192_mx0
      * conf_info_crt_lpi_1_dfm_167_160_mx0);
  assign nl_STORE_BATCH_LOOP_mul_1_nl = STORE_BATCH_LOOP_mul_2_nl * conf_info_crt_lpi_1_dfm_135_128_mx0;
  assign STORE_BATCH_LOOP_mul_1_nl = nl_STORE_BATCH_LOOP_mul_1_nl[15:0];
  assign STORE_BATCH_LOOP_mul_5_nl = conv_u2u_16_16(conf_info_crt_lpi_1_dfm_103_96_mx0
      * conf_info_crt_lpi_1_dfm_103_96_mx0);
  assign nl_STORE_BATCH_LOOP_mul_4_nl = STORE_BATCH_LOOP_mul_5_nl * conf_info_crt_lpi_1_dfm_135_128_mx0;
  assign STORE_BATCH_LOOP_mul_4_nl = nl_STORE_BATCH_LOOP_mul_4_nl[15:0];
  assign nl_STORE_BATCH_LOOP_mul_3_nl = STORE_BATCH_LOOP_mul_4_nl * conf_info_crt_lpi_1_dfm_71_64_mx0;
  assign STORE_BATCH_LOOP_mul_3_nl = nl_STORE_BATCH_LOOP_mul_3_nl[15:0];
  assign nl_STORE_BATCH_LOOP_acc_1_nl = STORE_BATCH_LOOP_mul_1_nl + STORE_BATCH_LOOP_mul_3_nl;
  assign STORE_BATCH_LOOP_acc_1_nl = nl_STORE_BATCH_LOOP_acc_1_nl[15:0];
  assign nl_STORE_BATCH_LOOP_mul_nl = STORE_BATCH_LOOP_acc_1_nl * conf_info_crt_lpi_1_dfm_231_224_mx0;
  assign STORE_BATCH_LOOP_mul_nl = nl_STORE_BATCH_LOOP_mul_nl[15:0];
  assign STORE_BATCH_LOOP_mul_8_nl = conv_u2u_16_16(n_w_out_lpi_1_dfm_3 * n_h_out_lpi_1_dfm_3);
  assign nl_STORE_BATCH_LOOP_mul_7_nl = STORE_BATCH_LOOP_mul_8_nl * conf_info_crt_lpi_1_dfm_135_128_mx0;
  assign STORE_BATCH_LOOP_mul_7_nl = nl_STORE_BATCH_LOOP_mul_7_nl[15:0];
  assign nl_STORE_BATCH_LOOP_mul_6_nl = STORE_BATCH_LOOP_mul_7_nl * STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1;
  assign STORE_BATCH_LOOP_mul_6_nl = nl_STORE_BATCH_LOOP_mul_6_nl[15:0];
  assign nl_dma_write_data_index_lpi_1_dfm_mx1w0 = STORE_BATCH_LOOP_mul_nl + STORE_BATCH_LOOP_mul_6_nl;
  assign dma_write_data_index_lpi_1_dfm_mx1w0 = nl_dma_write_data_index_lpi_1_dfm_mx1w0[15:0];
  assign conf_info_crt_lpi_1_dfm_199_192_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_199_192,
      (conf_info_rsci_idat_mxwt[55:48]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_167_160_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_167_160,
      (conf_info_rsci_idat_mxwt[47:40]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_135_128_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_135_128,
      (conf_info_rsci_idat_mxwt[39:32]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_103_96_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_103_96,
      (conf_info_rsci_idat_mxwt[31:24]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_71_64_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_71_64,
      (conf_info_rsci_idat_mxwt[23:16]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_231_224_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_231_224,
      (conf_info_rsci_idat_mxwt[63:56]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign operator_42_true_and_nl = (z_out_1[10]) & (z_out_1[0]);
  assign nl_operator_43_true_acc_nl = (z_out_1[8:1]) + conv_u2s_1_8(operator_42_true_and_nl)
      + 8'b00000001;
  assign operator_43_true_acc_nl = nl_operator_43_true_acc_nl[7:0];
  assign n_w_out_lpi_1_dfm_3 = MUX1HOT_v_8_3_2(n_w_out_lpi_1_dfm_1, (z_out_1[7:0]),
      operator_43_true_acc_nl, {(~ exitL_exit_STORE_BATCH_LOOP_sva) , STORE_BATCH_LOOP_asn_41
      , STORE_BATCH_LOOP_asn_43});
  assign operator_42_true_1_and_nl = (z_out[10]) & (z_out[0]);
  assign nl_operator_43_true_1_acc_nl = (z_out[8:1]) + conv_u2s_1_8(operator_42_true_1_and_nl)
      + 8'b00000001;
  assign operator_43_true_1_acc_nl = nl_operator_43_true_1_acc_nl[7:0];
  assign n_h_out_lpi_1_dfm_3 = MUX1HOT_v_8_3_2(n_h_out_lpi_1_dfm_1, (z_out[7:0]),
      operator_43_true_1_acc_nl, {(~ exitL_exit_STORE_BATCH_LOOP_sva) , STORE_BATCH_LOOP_asn_41
      , STORE_BATCH_LOOP_asn_43});
  assign exit_STORE_BATCH_LOOP_sva_2_mx0w0 = ~((~((STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1
      == (operator_8_false_4_acc_tmp[3:0])) & (operator_8_false_4_acc_tmp[7:4]==4'b0000)))
      | (operator_8_false_4_acc_tmp[8]));
  assign exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0 = ~(operator_8_false_2_acc_itm_4_1
      & or_139_cse);
  assign or_83_nl = or_dcpl_25 | and_dcpl_42;
  assign STORE_BATCH_LOOP_mux_8_nl = MUX_s_1_2_2(exit_STORE_BATCH_LOOP_sva_2_mx0w0,
      exit_STORE_BATCH_LOOP_sva_2, or_83_nl);
  assign exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0 = ((STORE_BATCH_LOOP_b_4_0_sva_2[4])
      | STORE_BATCH_LOOP_mux_8_nl) & exit_STORE_INNER_LOOP_lpi_1_dfm_3_mx0w0;
  assign STORE_INNER_LOOP_mux_1_nl = MUX_s_1_2_2(or_59_cse, exit_STORE_INNER_LOOP_lpi_1_dfm_1,
      or_dcpl_25);
  assign exit_STORE_INNER_LOOP_lpi_1_dfm_3_mx0w0 = STORE_INNER_LOOP_mux_1_nl & exit_STORE_INNER_LOOP_for_lpi_1_dfm_3_mx0w0;
  assign STORE_INNER_LOOP_for_mux_1_nl = MUX_s_1_2_2(exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0,
      exit_STORE_INNER_LOOP_for_lpi_1_dfm_1, and_162_cse);
  assign exit_STORE_INNER_LOOP_for_lpi_1_dfm_3_mx0w0 = STORE_INNER_LOOP_for_mux_1_nl
      & (~(operator_8_false_3_acc_itm_4_1 & or_138_cse));
  assign unequal_tmp_1 = ~((conf_info_rsci_idat_mxwt[7:0]==8'b00000001));
  assign operator_43_true_and_nl = (pad_acc_psp_sva_1[16]) & (pad_acc_psp_sva_1[0]);
  assign nl_operator_43_true_operator_43_true_acc_nl = (pad_acc_psp_sva_1[8:1]) +
      conv_u2s_1_8(operator_43_true_and_nl);
  assign operator_43_true_operator_43_true_acc_nl = nl_operator_43_true_operator_43_true_acc_nl[7:0];
  assign nl_pad_sva_1 = $signed(operator_43_true_operator_43_true_acc_nl) * $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[15:8]));
  assign pad_sva_1 = nl_pad_sva_1[7:0];
  assign nl_pad_acc_2_nl = ({1'b1 , (~ (conf_info_rsci_idat_mxwt[55:48]))}) + conv_u2s_8_9(conf_info_rsci_idat_mxwt[31:24])
      + 9'b000000001;
  assign pad_acc_2_nl = nl_pad_acc_2_nl[8:0];
  assign nl_operator_8_false_acc_nl = conv_u2s_8_9(conf_info_rsci_idat_mxwt[55:48])
      + 9'b111111111;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[8:0];
  assign nl_pad_mul_nl = $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[7:0])) * $signed(operator_8_false_acc_nl);
  assign pad_mul_nl = nl_pad_mul_nl[16:0];
  assign nl_pad_acc_psp_sva_1 = conv_s2s_9_17(pad_acc_2_nl) + pad_mul_nl;
  assign pad_acc_psp_sva_1 = nl_pad_acc_psp_sva_1[16:0];
  assign STORE_BATCH_LOOP_not_27_nl = ~ exitL_exit_STORE_BATCH_LOOP_sva;
  assign STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1 = MUX_v_4_2_2(4'b0000, STORE_BATCH_LOOP_b_4_0_lpi_1_3_0,
      STORE_BATCH_LOOP_not_27_nl);
  assign nl_STORE_BATCH_LOOP_b_4_0_sva_2 = conv_u2u_4_5(STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1)
      + 5'b00001;
  assign STORE_BATCH_LOOP_b_4_0_sva_2 = nl_STORE_BATCH_LOOP_b_4_0_sva_2[4:0];
  assign nl_operator_8_false_4_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_231_224_mx0)
      + 9'b111111111;
  assign operator_8_false_4_acc_tmp = nl_operator_8_false_4_acc_tmp[8:0];
  assign nl_STORE_INNER_LOOP_acc_tmp = conv_u2u_5_6(STORE_INNER_LOOP_fl_5_0_lpi_1_dfm_4_0_1)
      + 6'b000001;
  assign STORE_INNER_LOOP_acc_tmp = nl_STORE_INNER_LOOP_acc_tmp[5:0];
  assign STORE_INNER_LOOP_not_14_nl = ~ or_64_cse;
  assign STORE_INNER_LOOP_fl_5_0_lpi_1_dfm_4_0_1 = MUX_v_5_2_2(5'b00000, STORE_INNER_LOOP_fl_5_0_lpi_1_4_0,
      STORE_INNER_LOOP_not_14_nl);
  assign nl_operator_8_false_3_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_71_64_mx0)
      + 9'b111111111;
  assign operator_8_false_3_acc_tmp = nl_operator_8_false_3_acc_tmp[8:0];
  assign nl_operator_8_false_2_acc_nl = conv_u2s_4_5(STORE_INNER_LOOP_for_i_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_2_acc_nl = nl_operator_8_false_2_acc_nl[4:0];
  assign operator_8_false_2_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_2_acc_nl);
  assign nl_STORE_INNER_LOOP_for_i_4_0_sva_2 = STORE_INNER_LOOP_for_i_4_0_lpi_1_dfm_4
      + 5'b00001;
  assign STORE_INNER_LOOP_for_i_4_0_sva_2 = nl_STORE_INNER_LOOP_for_i_4_0_sva_2[4:0];
  assign STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_BATCH_LOOP_not_nl
      = ~ or_64_cse;
  assign STORE_INNER_LOOP_for_i_4_0_lpi_1_dfm_4 = MUX_v_5_2_2(5'b00000, STORE_INNER_LOOP_for_i_4_0_lpi_1,
      STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_BATCH_LOOP_not_nl);
  assign nl_operator_8_false_2_acc_tmp = conv_u2s_8_9(n_w_out_lpi_1_dfm_3) + 9'b111111111;
  assign operator_8_false_2_acc_tmp = nl_operator_8_false_2_acc_tmp[8:0];
  assign nl_operator_8_false_3_acc_nl = conv_u2s_4_5(STORE_INNER_LOOP_for_for_j_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_3_acc_nl = nl_operator_8_false_3_acc_nl[4:0];
  assign operator_8_false_3_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_3_acc_nl);
  assign nl_STORE_INNER_LOOP_for_for_j_4_0_sva_2 = STORE_INNER_LOOP_for_for_j_4_0_lpi_1_dfm_3
      + 5'b00001;
  assign STORE_INNER_LOOP_for_for_j_4_0_sva_2 = nl_STORE_INNER_LOOP_for_for_j_4_0_sva_2[4:0];
  assign STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_INNER_LOOP_nor_nl = ~(exit_STORE_INNER_LOOP_for_lpi_1_dfm_3
      | or_64_cse);
  assign STORE_INNER_LOOP_for_for_j_4_0_lpi_1_dfm_3 = MUX_v_5_2_2(5'b00000, STORE_INNER_LOOP_for_for_j_4_0_lpi_1,
      STORE_INNER_LOOP_STORE_INNER_LOOP_STORE_INNER_LOOP_nor_nl);
  assign STORE_INNER_LOOP_for_for_if_1_STORE_INNER_LOOP_for_for_if_1_nand_tmp = ~((STORE_INNER_LOOP_for_for_j_4_0_lpi_1_dfm_3
      == (operator_8_false_1_acc_tmp[4:0])) & (operator_8_false_1_acc_tmp[7:5]==3'b000));
  assign nl_operator_8_false_1_acc_tmp = conv_u2s_8_9(n_h_out_lpi_1_dfm_3) + 9'b111111111;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[8:0];
  assign main_stage_en_3 = or_5_cse & var_output_rsci_bawt & (dma_write_ctrl_rsci_bawt
      | (~ reg_dma_write_chnl_rsci_ivld_core_psct_cse)) & (dma_write_chnl_rsci_bawt
      | (~ reg_dma_write_chnl_rsci_ivld_core_psct_cse)) & (done_rsci_bawt | (~(exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2
      & main_stage_v_2)));
  assign STORE_BATCH_LOOP_asn_41 = (~ unequal_tmp_1) & exitL_exit_STORE_BATCH_LOOP_sva;
  assign STORE_BATCH_LOOP_asn_43 = unequal_tmp_1 & exitL_exit_STORE_BATCH_LOOP_sva;
  assign and_7_cse = exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2 & (~ done_rsci_bawt)
      & main_stage_v_2;
  assign or_tmp_7 = (~ main_stage_v_2) | done_rsci_bawt | (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2);
  assign and_165_cse = dma_write_chnl_rsci_bawt & dma_write_ctrl_rsci_bawt;
  assign and_tmp_4 = and_165_cse & or_tmp_7;
  assign mux_tmp_16 = MUX_s_1_2_2(or_tmp_7, and_tmp_4, reg_dma_write_chnl_rsci_ivld_core_psct_cse);
  assign and_tmp_5 = var_output_rsci_bawt & mux_tmp_16;
  assign nor_42_nl = ~(STORE_BATCH_LOOP_asn_itm | (~ and_tmp_5));
  assign mux_tmp_17 = MUX_s_1_2_2(nor_42_nl, and_tmp_5, conf_info_rsci_bawt);
  assign nand_tmp_4 = ~(exitL_exit_STORE_BATCH_LOOP_sva & (~ mux_tmp_17));
  assign or_tmp_40 = exitL_exit_STORE_BATCH_LOOP_sva | mux_tmp_17;
  assign nand_tmp_5 = ~(reg_dma_write_chnl_rsci_ivld_core_psct_cse & (~ and_165_cse));
  assign and_dcpl_9 = mux_tmp_16 & or_5_cse;
  assign and_dcpl_26 = exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2 & done_rsci_bawt &
      main_stage_v_2;
  assign and_dcpl_27 = (~(and_165_cse & reg_dma_write_chnl_rsci_ivld_core_psct_cse
      & exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1)) & and_dcpl_26;
  assign and_dcpl_28 = STORE_BATCH_LOOP_asn_itm & (~ conf_info_rsci_bawt);
  assign and_dcpl_30 = and_tmp_4 & (and_dcpl_28 | (~ var_output_rsci_bawt)) & reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  assign and_dcpl_34 = or_tmp_7 & reg_dma_write_chnl_rsci_ivld_core_psct_cse & dma_write_chnl_rsci_bawt
      & dma_write_ctrl_rsci_bawt;
  assign and_dcpl_42 = ~(nor_23_cse | (STORE_INNER_LOOP_acc_tmp[5]));
  assign and_dcpl_45 = (~ and_165_cse) & reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  assign or_dcpl_20 = and_7_cse | and_dcpl_45;
  assign or_dcpl_21 = or_dcpl_20 | and_dcpl_28;
  assign or_dcpl_22 = or_dcpl_21 | and_162_cse;
  assign or_dcpl_25 = and_162_cse | and_158_cse;
  assign or_89_nl = STORE_INNER_LOOP_for_for_if_1_STORE_INNER_LOOP_for_for_if_1_nand_tmp
      | (operator_8_false_1_acc_tmp[8]) | and_dcpl_45;
  assign mux_40_nl = MUX_s_1_2_2(and_dcpl_45, or_89_nl, operator_8_false_3_acc_itm_4_1);
  assign and_dcpl_46 = (~ mux_40_nl) & or_tmp_7;
  assign and_dcpl_53 = and_dcpl_46 & or_5_cse;
  assign and_dcpl_54 = and_dcpl_53 & exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0
      & var_output_rsci_bawt;
  assign and_dcpl_56 = mux_43_itm & or_tmp_7 & and_160_cse;
  assign or_dcpl_33 = ~(and_165_cse & reg_dma_write_chnl_rsci_ivld_core_psct_cse);
  assign mux_44_nl = MUX_s_1_2_2(nand_tmp_5, mux_43_itm, or_59_cse);
  assign mux_29_nl = MUX_s_1_2_2(nand_tmp_5, mux_44_nl, or_57_cse);
  assign mux_30_nl = MUX_s_1_2_2(nand_tmp_5, mux_29_nl, main_stage_en_3);
  assign or_tmp_56 = mux_30_nl & or_tmp_7 & var_output_rsci_bawt & STORE_BATCH_LOOP_asn_itm
      & conf_info_rsci_bawt & (fsm_output[1]);
  assign or_tmp_70 = mux_tmp_17 & (fsm_output[1]);
  assign main_stage_v_2_mx0c1 = ((~ exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2) | done_rsci_bawt)
      & main_stage_v_2 & or_dcpl_33;
  assign and_185_cse = ((conf_info_rsci_idat_mxwt[7:0]!=8'b00000001)) & (fsm_output[1]);
  assign if_if_and_cse = MUX_v_2_2_2(2'b00, (z_out_2[9:8]), and_185_cse);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (((~ mux_26_nl) & main_stage_en_3) | (fsm_output[0]) | or_tmp_56)
        ) begin
      reg_conf_info_rsci_iswt0_cse <= ~ or_tmp_56;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_var_output_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (main_stage_en_3 | (fsm_output[0])) ) begin
      reg_var_output_rsci_iswt0_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exitL_exit_STORE_BATCH_LOOP_sva <= 1'b1;
      dma_write_chnl_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2 <= 1'b0;
      exit_STORE_INNER_LOOP_lpi_1_dfm_3 <= 1'b0;
      exit_STORE_INNER_LOOP_for_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( STORE_BATCH_LOOP_and_2_cse ) begin
      exitL_exit_STORE_BATCH_LOOP_sva <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
      dma_write_chnl_rsci_idat_31_0 <= var_output_rsci_idat_mxwt;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
      exit_STORE_INNER_LOOP_lpi_1_dfm_3 <= exit_STORE_INNER_LOOP_lpi_1_dfm_3_mx0w0;
      exit_STORE_INNER_LOOP_for_lpi_1_dfm_3 <= exit_STORE_INNER_LOOP_for_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_rsci_idat_15_0 <= 16'b0000000000000000;
    end
    else if ( core_wen & (~ (fsm_output[0])) & ((and_dcpl_9 & or_64_cse & var_output_rsci_bawt)
        | and_34_rgt) ) begin
      dma_write_ctrl_rsci_idat_15_0 <= MUX_v_16_2_2(dma_write_data_index_lpi_1_dfm_mx1w0,
          dma_write_data_index_lpi_1, and_34_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_done_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((or_tmp_7 & dma_write_ctrl_rsci_bawt & dma_write_chnl_rsci_bawt
        & reg_dma_write_chnl_rsci_ivld_core_psct_cse & exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1)
        | and_dcpl_27) ) begin
      reg_done_rsci_ivld_core_psct_cse <= ~ and_dcpl_27;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_write_chnl_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_70 | and_dcpl_30) ) begin
      reg_dma_write_chnl_rsci_ivld_core_psct_cse <= ~ and_dcpl_30;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_asn_itm <= 1'b1;
    end
    else if ( core_wen & ((main_stage_en_3 & (fsm_output[1])) | ((~ STORE_BATCH_LOOP_asn_itm)
        & main_stage_en_3)) ) begin
      STORE_BATCH_LOOP_asn_itm <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_crt_lpi_1_dfm_199_192 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_167_160 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_135_128 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_103_96 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_71_64 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_231_224 <= 8'b00000000;
    end
    else if ( core_wen ) begin
      conf_info_crt_lpi_1_dfm_199_192 <= conf_info_crt_lpi_1_dfm_199_192_mx0;
      conf_info_crt_lpi_1_dfm_167_160 <= conf_info_crt_lpi_1_dfm_167_160_mx0;
      conf_info_crt_lpi_1_dfm_135_128 <= conf_info_crt_lpi_1_dfm_135_128_mx0;
      conf_info_crt_lpi_1_dfm_103_96 <= conf_info_crt_lpi_1_dfm_103_96_mx0;
      conf_info_crt_lpi_1_dfm_71_64 <= conf_info_crt_lpi_1_dfm_71_64_mx0;
      conf_info_crt_lpi_1_dfm_231_224 <= conf_info_crt_lpi_1_dfm_231_224_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      n_w_out_lpi_1_dfm_1 <= 8'b00000000;
      n_h_out_lpi_1_dfm_1 <= 8'b00000000;
      dma_write_data_index_lpi_1 <= 16'b0000000000000000;
    end
    else if ( n_w_out_and_cse ) begin
      n_w_out_lpi_1_dfm_1 <= n_w_out_lpi_1_dfm_3;
      n_h_out_lpi_1_dfm_1 <= n_h_out_lpi_1_dfm_3;
      dma_write_data_index_lpi_1 <= nl_dma_write_data_index_lpi_1[15:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_22 | and_158_cse | and_dcpl_42 | (~ var_output_rsci_bawt)
        | (fsm_output[0]))) ) begin
      exit_STORE_BATCH_LOOP_sva_2 <= exit_STORE_BATCH_LOOP_sva_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_INNER_LOOP_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_22 | and_158_cse | (~ var_output_rsci_bawt) |
        (fsm_output[0]))) ) begin
      exit_STORE_INNER_LOOP_lpi_1_dfm_1 <= or_59_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_INNER_LOOP_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_21 | and_162_cse | (~ var_output_rsci_bawt) |
        (fsm_output[0]))) ) begin
      exit_STORE_INNER_LOOP_for_lpi_1_dfm_1 <= exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_INNER_LOOP_for_for_j_4_0_lpi_1 <= 5'b00000;
    end
    else if ( core_wen & ((and_dcpl_46 & and_160_cse) | and_64_rgt) ) begin
      STORE_INNER_LOOP_for_for_j_4_0_lpi_1 <= MUX_v_5_2_2(({{4{exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0}},
          exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0}), STORE_INNER_LOOP_for_for_j_4_0_sva_2,
          and_64_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_INNER_LOOP_for_i_4_0_lpi_1 <= 5'b00000;
    end
    else if ( core_wen & (and_dcpl_54 | STORE_INNER_LOOP_for_and_3_rgt | STORE_INNER_LOOP_for_and_4_rgt)
        ) begin
      STORE_INNER_LOOP_for_i_4_0_lpi_1 <= MUX1HOT_v_5_3_2(({{4{or_59_cse}}, or_59_cse}),
          STORE_INNER_LOOP_for_i_4_0_sva_2, STORE_INNER_LOOP_for_i_4_0_lpi_1_dfm_4,
          {and_dcpl_54 , STORE_INNER_LOOP_for_and_3_rgt , STORE_INNER_LOOP_for_and_4_rgt});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_INNER_LOOP_fl_5_0_lpi_1_4_0 <= 5'b00000;
    end
    else if ( core_wen & (and_dcpl_54 | and_dcpl_56) ) begin
      STORE_INNER_LOOP_fl_5_0_lpi_1_4_0 <= MUX_v_5_2_2((STORE_INNER_LOOP_acc_tmp[4:0]),
          STORE_INNER_LOOP_fl_5_0_lpi_1_dfm_4_0_1, and_dcpl_56);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_b_4_0_lpi_1_3_0 <= 4'b0000;
    end
    else if ( core_wen & ((and_dcpl_53 & exit_STORE_INNER_LOOP_for_lpi_1_dfm_1_mx0w0
        & or_59_cse & var_output_rsci_bawt) | and_76_rgt) ) begin
      STORE_BATCH_LOOP_b_4_0_lpi_1_3_0 <= MUX_v_4_2_2((STORE_BATCH_LOOP_b_4_0_sva_2[3:0]),
          STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1, and_76_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_20) ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_34 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2 <= 1'b0;
    end
    else if ( core_wen & (~(and_7_cse | or_dcpl_33)) ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1;
    end
  end
  assign mux_22_nl = MUX_s_1_2_2((~ or_tmp_40), nand_tmp_4, or_138_cse);
  assign mux_23_nl = MUX_s_1_2_2((~ or_tmp_40), mux_22_nl, operator_8_false_3_acc_itm_4_1);
  assign mux_24_nl = MUX_s_1_2_2(mux_23_nl, nand_tmp_4, and_158_cse);
  assign mux_25_nl = MUX_s_1_2_2(nand_tmp_4, mux_24_nl, or_59_cse);
  assign mux_26_nl = MUX_s_1_2_2(nand_tmp_4, mux_25_nl, or_57_cse);
  assign nor_41_nl = ~(exitL_exit_STORE_BATCH_LOOP_sva | exit_STORE_INNER_LOOP_lpi_1_dfm_3
      | exit_STORE_BATCH_LOOP_lpi_1_dfm_2);
  assign dma_write_data_index_mux_1_nl = MUX_v_16_2_2(dma_write_data_index_lpi_1_dfm_mx1w0,
      dma_write_data_index_lpi_1, nor_41_nl);
  assign nl_dma_write_data_index_lpi_1  = dma_write_data_index_mux_1_nl + 16'b0000000000000001;
  assign if_if_nand_2_cse = ~(and_185_cse & (~((conf_info_rsci_idat_mxwt[7:0]==8'b00000001)
      & (fsm_output[1]))));
  assign nl_acc_nl = conv_u2u_11_12({if_if_and_cse , (z_out_2[7:0]) , if_if_nand_2_cse})
      + conv_s2u_10_12({and_185_cse , (conf_info_rsci_idat_mxwt[47:40]) , 1'b1});
  assign acc_nl = nl_acc_nl[11:0];
  assign z_out = readslicef_12_11_1(acc_nl);
  assign nl_acc_1_nl = conv_u2u_11_12({if_if_and_cse , (z_out_2[7:0]) , if_if_nand_2_cse})
      + conv_s2u_10_12({and_185_cse , (conf_info_rsci_idat_mxwt[55:48]) , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[11:0];
  assign z_out_1 = readslicef_12_11_1(acc_1_nl);
  assign if_if_and_3_nl = (pad_sva_1[7]) & and_185_cse;
  assign nl_acc_2_nl = conv_u2u_10_11({if_if_and_3_nl , (pad_sva_1[6:0]) , 2'b01})
      + conv_u2u_9_11({(~ (conf_info_rsci_idat_mxwt[31:24])) , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[10:0];
  assign z_out_2 = readslicef_11_10_1(acc_2_nl);

  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [16:0] conv_s2s_9_17 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_17 = {{8{vector[8]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_10_12 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_12 = {{2{vector[9]}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_16 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core (
  clk, rst, acc_done_rsc_vld, config_done_cns_rdy, config_done_cns_vld, load_done_cns_rdy,
      load_done_cns_vld, compute_done_cns_rdy, compute_done_cns_vld, store_done_cns_rdy,
      store_done_cns_vld
);
  input clk;
  input rst;
  output acc_done_rsc_vld;
  output config_done_cns_rdy;
  input config_done_cns_vld;
  output load_done_cns_rdy;
  input load_done_cns_vld;
  output compute_done_cns_rdy;
  input compute_done_cns_vld;
  output store_done_cns_rdy;
  input store_done_cns_vld;



  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core_core conv2dlb_cxx_catapult_core_core_inst
      (
      .clk(clk),
      .rst(rst),
      .acc_done_rsc_vld(acc_done_rsc_vld),
      .config_done_cns_rdy(config_done_cns_rdy),
      .config_done_cns_vld(config_done_cns_vld),
      .load_done_cns_rdy(load_done_cns_rdy),
      .load_done_cns_vld(load_done_cns_vld),
      .compute_done_cns_rdy(compute_done_cns_rdy),
      .compute_done_cns_vld(compute_done_cns_vld),
      .store_done_cns_rdy(store_done_cns_rdy),
      .store_done_cns_vld(store_done_cns_vld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_config
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_config (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_conf_load_rsc_dat,
      plm_conf_load_rsc_vld, plm_conf_load_rsc_rdy, plm_conf_compute_rsc_dat, plm_conf_compute_rsc_vld,
      plm_conf_compute_rsc_rdy, plm_conf_store_rsc_dat, plm_conf_store_rsc_vld, plm_conf_store_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [255:0] plm_conf_load_rsc_dat;
  output plm_conf_load_rsc_vld;
  input plm_conf_load_rsc_rdy;
  output [255:0] plm_conf_compute_rsc_dat;
  output plm_conf_compute_rsc_vld;
  input plm_conf_compute_rsc_rdy;
  output [255:0] plm_conf_store_rsc_dat;
  output plm_conf_store_rsc_vld;
  input plm_conf_store_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;



  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_config_core config_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .plm_conf_load_rsc_dat(plm_conf_load_rsc_dat),
      .plm_conf_load_rsc_vld(plm_conf_load_rsc_vld),
      .plm_conf_load_rsc_rdy(plm_conf_load_rsc_rdy),
      .plm_conf_compute_rsc_dat(plm_conf_compute_rsc_dat),
      .plm_conf_compute_rsc_vld(plm_conf_compute_rsc_vld),
      .plm_conf_compute_rsc_rdy(plm_conf_compute_rsc_rdy),
      .plm_conf_store_rsc_dat(plm_conf_store_rsc_dat),
      .plm_conf_store_rsc_vld(plm_conf_store_rsc_vld),
      .plm_conf_store_rsc_rdy(plm_conf_store_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_load
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_load (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, buf_linear_rsc_dat,
      buf_linear_rsc_vld, buf_linear_rsc_rdy, plm_kernel_rsc_dat, plm_kernel_rsc_vld,
      plm_kernel_rsc_rdy, dma_read_ctrl_rsc_dat, dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy,
      dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy, done_rsc_rdy,
      done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [4031:0] buf_linear_rsc_dat;
  output buf_linear_rsc_vld;
  input buf_linear_rsc_rdy;
  output [1567:0] plm_kernel_rsc_dat;
  output plm_kernel_rsc_vld;
  input plm_kernel_rsc_rdy;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d;
  wire [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d;
  wire [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d;
  wire [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_clken;
  wire [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_q;
  wire [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_radr;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_we;
  wire [31:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_d;
  wire [13:0] LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wadr;
  wire LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd14),
  .data_width(32'sd32),
  .depth(32'sd10368),
  .latency(32'sd1)) LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_comp (
      .clk(clk),
      .clken(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_clken),
      .d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_d),
      .q(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_q),
      .radr(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_radr),
      .wadr(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wadr),
      .we(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_we)
    );
  esp_acc_conv2dlb_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_12_14_32_10368_10368_32_1_gen
      LOAD_BATCH_LOOP_plm_tmp_in_data_rsci (
      .clken(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_clken),
      .q(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_q),
      .radr(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_radr),
      .we(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_we),
      .d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_d),
      .wadr(LOAD_BATCH_LOOP_plm_tmp_in_data_rsc_wadr),
      .clken_d(1'b1),
      .d_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d),
      .q_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d),
      .radr_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d),
      .wadr_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d),
      .we_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_conv2dlb_cxx_catapult_load_core load_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .buf_linear_rsc_dat(buf_linear_rsc_dat),
      .buf_linear_rsc_vld(buf_linear_rsc_vld),
      .buf_linear_rsc_rdy(buf_linear_rsc_rdy),
      .plm_kernel_rsc_dat(plm_kernel_rsc_dat),
      .plm_kernel_rsc_vld(plm_kernel_rsc_vld),
      .plm_kernel_rsc_rdy(plm_kernel_rsc_rdy),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_d_d),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_q_d),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_radr_d),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_wadr_d),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_pff(LOAD_BATCH_LOOP_plm_tmp_in_data_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_compute
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_compute (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, buf_linear_rsc_dat,
      buf_linear_rsc_vld, buf_linear_rsc_rdy, plm_kernel_rsc_dat, plm_kernel_rsc_vld,
      plm_kernel_rsc_rdy, var_output_rsc_dat, var_output_rsc_vld, var_output_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input [4031:0] buf_linear_rsc_dat;
  input buf_linear_rsc_vld;
  output buf_linear_rsc_rdy;
  input [1567:0] plm_kernel_rsc_dat;
  input plm_kernel_rsc_vld;
  output plm_kernel_rsc_rdy;
  output [31:0] var_output_rsc_dat;
  output var_output_rsc_vld;
  input var_output_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;



  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_compute_core compute_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .buf_linear_rsc_dat(buf_linear_rsc_dat),
      .buf_linear_rsc_vld(buf_linear_rsc_vld),
      .buf_linear_rsc_rdy(buf_linear_rsc_rdy),
      .plm_kernel_rsc_dat(plm_kernel_rsc_dat),
      .plm_kernel_rsc_vld(plm_kernel_rsc_vld),
      .plm_kernel_rsc_rdy(plm_kernel_rsc_rdy),
      .var_output_rsc_dat(var_output_rsc_dat),
      .var_output_rsc_vld(var_output_rsc_vld),
      .var_output_rsc_rdy(var_output_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_store
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_store (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, var_output_rsc_dat,
      var_output_rsc_vld, var_output_rsc_rdy, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld,
      dma_write_ctrl_rsc_rdy, dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input [31:0] var_output_rsc_dat;
  input var_output_rsc_vld;
  output var_output_rsc_rdy;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;



  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2dlb_cxx_catapult_store_core store_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .var_output_rsc_dat(var_output_rsc_dat),
      .var_output_rsc_vld(var_output_rsc_vld),
      .var_output_rsc_rdy(var_output_rsc_rdy),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_struct
// ------------------------------------------------------------------


module esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_struct (
  clk, rst, conf_info_rsc_dat_batch, conf_info_rsc_dat_n_w, conf_info_rsc_dat_n_h,
      conf_info_rsc_dat_n_c, conf_info_rsc_dat_kern, conf_info_rsc_dat_filt, conf_info_rsc_dat_same,
      conf_info_rsc_dat_stride, conf_info_rsc_vld, conf_info_rsc_rdy, dma_read_ctrl_rsc_dat_size,
      dma_read_ctrl_rsc_dat_length, dma_read_ctrl_rsc_dat_index, dma_read_ctrl_rsc_vld,
      dma_read_ctrl_rsc_rdy, dma_write_ctrl_rsc_dat_size, dma_write_ctrl_rsc_dat_length,
      dma_write_ctrl_rsc_dat_index, dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy,
      dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy, dma_write_chnl_rsc_dat,
      dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, acc_done_rsc_vld
);
  input clk;
  input rst;
  input [31:0] conf_info_rsc_dat_batch;
  input [31:0] conf_info_rsc_dat_n_w;
  input [31:0] conf_info_rsc_dat_n_h;
  input [31:0] conf_info_rsc_dat_n_c;
  input [31:0] conf_info_rsc_dat_kern;
  input [31:0] conf_info_rsc_dat_filt;
  input [31:0] conf_info_rsc_dat_same;
  input [31:0] conf_info_rsc_dat_stride;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [2:0] dma_read_ctrl_rsc_dat_size;
  output [31:0] dma_read_ctrl_rsc_dat_length;
  output [31:0] dma_read_ctrl_rsc_dat_index;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  output [2:0] dma_write_ctrl_rsc_dat_size;
  output [31:0] dma_write_ctrl_rsc_dat_length;
  output [31:0] dma_write_ctrl_rsc_dat_index;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  output acc_done_rsc_vld;


  // Interconnect Declarations
  wire [255:0] plm_conf_load_rsc_dat_nconfig_inst;
  wire plm_conf_load_rsc_rdy_nconfig_inst;
  wire [255:0] plm_conf_compute_rsc_dat_nconfig_inst;
  wire plm_conf_compute_rsc_rdy_nconfig_inst;
  wire [255:0] plm_conf_store_rsc_dat_nconfig_inst;
  wire plm_conf_store_rsc_rdy_nconfig_inst;
  wire done_rsc_rdy_nconfig_inst;
  wire [255:0] conf_info_rsc_dat_nload_inst;
  wire conf_info_rsc_vld_nload_inst;
  wire [4031:0] buf_linear_rsc_dat_nload_inst;
  wire buf_linear_rsc_rdy_nload_inst;
  wire [1567:0] plm_kernel_rsc_dat_nload_inst;
  wire plm_kernel_rsc_rdy_nload_inst;
  wire [66:0] dma_read_ctrl_rsc_dat_nload_inst;
  wire done_rsc_rdy_nload_inst;
  wire [255:0] conf_info_rsc_dat_ncompute_inst;
  wire conf_info_rsc_vld_ncompute_inst;
  wire [4031:0] buf_linear_rsc_dat_ncompute_inst;
  wire buf_linear_rsc_vld_ncompute_inst;
  wire [1567:0] plm_kernel_rsc_dat_ncompute_inst;
  wire plm_kernel_rsc_vld_ncompute_inst;
  wire [31:0] var_output_rsc_dat_ncompute_inst;
  wire var_output_rsc_rdy_ncompute_inst;
  wire done_rsc_rdy_ncompute_inst;
  wire [255:0] conf_info_rsc_dat_nstore_inst;
  wire conf_info_rsc_vld_nstore_inst;
  wire [31:0] var_output_rsc_dat_nstore_inst;
  wire var_output_rsc_vld_nstore_inst;
  wire [66:0] dma_write_ctrl_rsc_dat_nstore_inst;
  wire [63:0] dma_write_chnl_rsc_dat_nstore_inst;
  wire done_rsc_rdy_nstore_inst;
  wire config_done_cns_vld_nconv2dlb_cxx_catapult_core_inst;
  wire load_done_cns_vld_nconv2dlb_cxx_catapult_core_inst;
  wire compute_done_cns_vld_nconv2dlb_cxx_catapult_core_inst;
  wire store_done_cns_vld_nconv2dlb_cxx_catapult_core_inst;
  wire conf_info_rsc_rdy_nconfig_inst_bud;
  wire plm_conf_load_rsc_vld_nconfig_inst_bud;
  wire conf_info_rsc_rdy_nload_inst_bud;
  wire plm_conf_compute_rsc_vld_nconfig_inst_bud;
  wire conf_info_rsc_rdy_ncompute_inst_bud;
  wire plm_conf_store_rsc_vld_nconfig_inst_bud;
  wire conf_info_rsc_rdy_nstore_inst_bud;
  wire done_rsc_vld_nconfig_inst_bud;
  wire config_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud;
  wire buf_linear_rsc_vld_nload_inst_bud;
  wire buf_linear_rsc_rdy_ncompute_inst_bud;
  wire plm_kernel_rsc_vld_nload_inst_bud;
  wire plm_kernel_rsc_rdy_ncompute_inst_bud;
  wire dma_read_ctrl_rsc_vld_nload_inst_bud;
  wire dma_read_chnl_rsc_rdy_nload_inst_bud;
  wire done_rsc_vld_nload_inst_bud;
  wire load_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud;
  wire var_output_rsc_vld_ncompute_inst_bud;
  wire var_output_rsc_rdy_nstore_inst_bud;
  wire done_rsc_vld_ncompute_inst_bud;
  wire compute_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud;
  wire dma_write_ctrl_rsc_vld_nstore_inst_bud;
  wire dma_write_chnl_rsc_vld_nstore_inst_bud;
  wire done_rsc_vld_nstore_inst_bud;
  wire store_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud;
  wire acc_done_rsc_vld_nconv2dlb_cxx_catapult_core_inst_bud;
  wire plm_conf_load_unc_2;
  wire plm_conf_load_idle;
  wire plm_conf_compute_unc_2;
  wire plm_conf_compute_idle;
  wire plm_conf_store_unc_2;
  wire plm_conf_store_idle;
  wire buf_linear_unc_2;
  wire buf_linear_idle;
  wire plm_kernel_unc_2;
  wire plm_kernel_idle;
  wire var_output_unc_2;
  wire var_output_idle;


  // Interconnect Declarations for Component Instantiations 
  wire [255:0] nl_config_inst_conf_info_rsc_dat;
  assign nl_config_inst_conf_info_rsc_dat = {conf_info_rsc_dat_batch , conf_info_rsc_dat_n_w
      , conf_info_rsc_dat_n_h , conf_info_rsc_dat_n_c , conf_info_rsc_dat_kern ,
      conf_info_rsc_dat_filt , conf_info_rsc_dat_same , conf_info_rsc_dat_stride};
  esp_acc_conv2dlb_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd37),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_conf_load_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_conf_load_rsc_rdy_nconfig_inst),
      .din_vld(plm_conf_load_rsc_vld_nconfig_inst_bud),
      .din(plm_conf_load_rsc_dat_nconfig_inst),
      .dout_rdy(conf_info_rsc_rdy_nload_inst_bud),
      .dout_vld(conf_info_rsc_vld_nload_inst),
      .dout(conf_info_rsc_dat_nload_inst),
      .sz(plm_conf_load_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_conf_load_idle)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd38),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_conf_compute_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_conf_compute_rsc_rdy_nconfig_inst),
      .din_vld(plm_conf_compute_rsc_vld_nconfig_inst_bud),
      .din(plm_conf_compute_rsc_dat_nconfig_inst),
      .dout_rdy(conf_info_rsc_rdy_ncompute_inst_bud),
      .dout_vld(conf_info_rsc_vld_ncompute_inst),
      .dout(conf_info_rsc_dat_ncompute_inst),
      .sz(plm_conf_compute_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_conf_compute_idle)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd39),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_conf_store_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_conf_store_rsc_rdy_nconfig_inst),
      .din_vld(plm_conf_store_rsc_vld_nconfig_inst_bud),
      .din(plm_conf_store_rsc_dat_nconfig_inst),
      .dout_rdy(conf_info_rsc_rdy_nstore_inst_bud),
      .dout_vld(conf_info_rsc_vld_nstore_inst),
      .dout(conf_info_rsc_dat_nstore_inst),
      .sz(plm_conf_store_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_conf_store_idle)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd40)) config_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_nconfig_inst_bud),
      .dout_vld(done_rsc_rdy_nconfig_inst),
      .din_vld(config_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .din_rdy(config_done_cns_vld_nconv2dlb_cxx_catapult_core_inst)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd34),
  .width(32'sd4032),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) buf_linear_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(buf_linear_rsc_rdy_nload_inst),
      .din_vld(buf_linear_rsc_vld_nload_inst_bud),
      .din(buf_linear_rsc_dat_nload_inst),
      .dout_rdy(buf_linear_rsc_rdy_ncompute_inst_bud),
      .dout_vld(buf_linear_rsc_vld_ncompute_inst),
      .dout(buf_linear_rsc_dat_ncompute_inst),
      .sz(buf_linear_unc_2),
      .sz_req(1'b0),
      .is_idle(buf_linear_idle)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd35),
  .width(32'sd1568),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_kernel_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_kernel_rsc_rdy_nload_inst),
      .din_vld(plm_kernel_rsc_vld_nload_inst_bud),
      .din(plm_kernel_rsc_dat_nload_inst),
      .dout_rdy(plm_kernel_rsc_rdy_ncompute_inst_bud),
      .dout_vld(plm_kernel_rsc_vld_ncompute_inst),
      .dout(plm_kernel_rsc_dat_ncompute_inst),
      .sz(plm_kernel_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_kernel_idle)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd41)) load_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_nload_inst_bud),
      .dout_vld(done_rsc_rdy_nload_inst),
      .din_vld(load_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .din_rdy(load_done_cns_vld_nconv2dlb_cxx_catapult_core_inst)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd36),
  .width(32'sd32),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) var_output_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(var_output_rsc_rdy_ncompute_inst),
      .din_vld(var_output_rsc_vld_ncompute_inst_bud),
      .din(var_output_rsc_dat_ncompute_inst),
      .dout_rdy(var_output_rsc_rdy_nstore_inst_bud),
      .dout_vld(var_output_rsc_vld_nstore_inst),
      .dout(var_output_rsc_dat_nstore_inst),
      .sz(var_output_unc_2),
      .sz_req(1'b0),
      .is_idle(var_output_idle)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd42)) compute_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_ncompute_inst_bud),
      .dout_vld(done_rsc_rdy_ncompute_inst),
      .din_vld(compute_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .din_rdy(compute_done_cns_vld_nconv2dlb_cxx_catapult_core_inst)
    );
  esp_acc_conv2dlb_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd43)) store_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_nstore_inst_bud),
      .dout_vld(done_rsc_rdy_nstore_inst),
      .din_vld(store_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .din_rdy(store_done_cns_vld_nconv2dlb_cxx_catapult_core_inst)
    );
  esp_acc_conv2dlb_cxx_catapult_config config_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(nl_config_inst_conf_info_rsc_dat[255:0]),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_nconfig_inst_bud),
      .plm_conf_load_rsc_dat(plm_conf_load_rsc_dat_nconfig_inst),
      .plm_conf_load_rsc_vld(plm_conf_load_rsc_vld_nconfig_inst_bud),
      .plm_conf_load_rsc_rdy(plm_conf_load_rsc_rdy_nconfig_inst),
      .plm_conf_compute_rsc_dat(plm_conf_compute_rsc_dat_nconfig_inst),
      .plm_conf_compute_rsc_vld(plm_conf_compute_rsc_vld_nconfig_inst_bud),
      .plm_conf_compute_rsc_rdy(plm_conf_compute_rsc_rdy_nconfig_inst),
      .plm_conf_store_rsc_dat(plm_conf_store_rsc_dat_nconfig_inst),
      .plm_conf_store_rsc_vld(plm_conf_store_rsc_vld_nconfig_inst_bud),
      .plm_conf_store_rsc_rdy(plm_conf_store_rsc_rdy_nconfig_inst),
      .done_rsc_rdy(done_rsc_rdy_nconfig_inst),
      .done_rsc_vld(done_rsc_vld_nconfig_inst_bud)
    );
  esp_acc_conv2dlb_cxx_catapult_load load_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat_nload_inst),
      .conf_info_rsc_vld(conf_info_rsc_vld_nload_inst),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_nload_inst_bud),
      .buf_linear_rsc_dat(buf_linear_rsc_dat_nload_inst),
      .buf_linear_rsc_vld(buf_linear_rsc_vld_nload_inst_bud),
      .buf_linear_rsc_rdy(buf_linear_rsc_rdy_nload_inst),
      .plm_kernel_rsc_dat(plm_kernel_rsc_dat_nload_inst),
      .plm_kernel_rsc_vld(plm_kernel_rsc_vld_nload_inst_bud),
      .plm_kernel_rsc_rdy(plm_kernel_rsc_rdy_nload_inst),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat_nload_inst),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld_nload_inst_bud),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy_nload_inst_bud),
      .done_rsc_rdy(done_rsc_rdy_nload_inst),
      .done_rsc_vld(done_rsc_vld_nload_inst_bud)
    );
  esp_acc_conv2dlb_cxx_catapult_compute compute_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat_ncompute_inst),
      .conf_info_rsc_vld(conf_info_rsc_vld_ncompute_inst),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_ncompute_inst_bud),
      .buf_linear_rsc_dat(buf_linear_rsc_dat_ncompute_inst),
      .buf_linear_rsc_vld(buf_linear_rsc_vld_ncompute_inst),
      .buf_linear_rsc_rdy(buf_linear_rsc_rdy_ncompute_inst_bud),
      .plm_kernel_rsc_dat(plm_kernel_rsc_dat_ncompute_inst),
      .plm_kernel_rsc_vld(plm_kernel_rsc_vld_ncompute_inst),
      .plm_kernel_rsc_rdy(plm_kernel_rsc_rdy_ncompute_inst_bud),
      .var_output_rsc_dat(var_output_rsc_dat_ncompute_inst),
      .var_output_rsc_vld(var_output_rsc_vld_ncompute_inst_bud),
      .var_output_rsc_rdy(var_output_rsc_rdy_ncompute_inst),
      .done_rsc_rdy(done_rsc_rdy_ncompute_inst),
      .done_rsc_vld(done_rsc_vld_ncompute_inst_bud)
    );
  esp_acc_conv2dlb_cxx_catapult_store store_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat_nstore_inst),
      .conf_info_rsc_vld(conf_info_rsc_vld_nstore_inst),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_nstore_inst_bud),
      .var_output_rsc_dat(var_output_rsc_dat_nstore_inst),
      .var_output_rsc_vld(var_output_rsc_vld_nstore_inst),
      .var_output_rsc_rdy(var_output_rsc_rdy_nstore_inst_bud),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat_nstore_inst),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld_nstore_inst_bud),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat_nstore_inst),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld_nstore_inst_bud),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy_nstore_inst),
      .done_rsc_vld(done_rsc_vld_nstore_inst_bud)
    );
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_core conv2dlb_cxx_catapult_core_inst
      (
      .clk(clk),
      .rst(rst),
      .acc_done_rsc_vld(acc_done_rsc_vld_nconv2dlb_cxx_catapult_core_inst_bud),
      .config_done_cns_rdy(config_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .config_done_cns_vld(config_done_cns_vld_nconv2dlb_cxx_catapult_core_inst),
      .load_done_cns_rdy(load_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .load_done_cns_vld(load_done_cns_vld_nconv2dlb_cxx_catapult_core_inst),
      .compute_done_cns_rdy(compute_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .compute_done_cns_vld(compute_done_cns_vld_nconv2dlb_cxx_catapult_core_inst),
      .store_done_cns_rdy(store_done_cns_rdy_nconv2dlb_cxx_catapult_core_inst_bud),
      .store_done_cns_vld(store_done_cns_vld_nconv2dlb_cxx_catapult_core_inst)
    );
  assign conf_info_rsc_rdy = conf_info_rsc_rdy_nconfig_inst_bud;
  assign dma_read_ctrl_rsc_dat_index = dma_read_ctrl_rsc_dat_nload_inst[31:0];
  assign dma_read_ctrl_rsc_dat_length = dma_read_ctrl_rsc_dat_nload_inst[63:32];
  assign dma_read_ctrl_rsc_dat_size = dma_read_ctrl_rsc_dat_nload_inst[66:64];
  assign dma_write_ctrl_rsc_dat_index = dma_write_ctrl_rsc_dat_nstore_inst[31:0];
  assign dma_write_ctrl_rsc_dat_length = dma_write_ctrl_rsc_dat_nstore_inst[63:32];
  assign dma_write_ctrl_rsc_dat_size = dma_write_ctrl_rsc_dat_nstore_inst[66:64];
  assign dma_read_ctrl_rsc_vld = dma_read_ctrl_rsc_vld_nload_inst_bud;
  assign dma_read_chnl_rsc_rdy = dma_read_chnl_rsc_rdy_nload_inst_bud;
  assign dma_write_ctrl_rsc_vld = dma_write_ctrl_rsc_vld_nstore_inst_bud;
  assign dma_write_chnl_rsc_vld = dma_write_chnl_rsc_vld_nstore_inst_bud;
  assign dma_write_chnl_rsc_dat = dma_write_chnl_rsc_dat_nstore_inst;
  assign acc_done_rsc_vld = acc_done_rsc_vld_nconv2dlb_cxx_catapult_core_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv2dlb_cxx_catapult_hier_fx32_dma64
// ------------------------------------------------------------------


module conv2dlb_cxx_catapult_hier_fx32_dma64 (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, dma_read_ctrl_rsc_dat,
      dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld,
      dma_write_ctrl_rsc_rdy, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy,
      dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, acc_done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  output acc_done_rsc_vld;


  // Interconnect Declarations
  wire [2:0] dma_read_ctrl_rsc_dat_size;
  wire [31:0] dma_read_ctrl_rsc_dat_length;
  wire [31:0] dma_read_ctrl_rsc_dat_index;
  wire [2:0] dma_write_ctrl_rsc_dat_size;
  wire [31:0] dma_write_ctrl_rsc_dat_length;
  wire [31:0] dma_write_ctrl_rsc_dat_index;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_batch;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_batch = conf_info_rsc_dat[255:224];
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w = conf_info_rsc_dat[223:192];
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h = conf_info_rsc_dat[191:160];
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c = conf_info_rsc_dat[159:128];
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_kern;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_kern = conf_info_rsc_dat[127:96];
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_filt;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_filt = conf_info_rsc_dat[95:64];
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_same;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_same = conf_info_rsc_dat[63:32];
  wire [31:0] nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_stride;
  assign nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_stride = conf_info_rsc_dat[31:0];
  esp_acc_conv2dlb_cxx_catapult_conv2dlb_cxx_catapult_struct conv2dlb_cxx_catapult_struct_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat_batch(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_batch[31:0]),
      .conf_info_rsc_dat_n_w(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w[31:0]),
      .conf_info_rsc_dat_n_h(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h[31:0]),
      .conf_info_rsc_dat_n_c(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c[31:0]),
      .conf_info_rsc_dat_kern(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_kern[31:0]),
      .conf_info_rsc_dat_filt(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_filt[31:0]),
      .conf_info_rsc_dat_same(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_same[31:0]),
      .conf_info_rsc_dat_stride(nl_conv2dlb_cxx_catapult_struct_inst_conf_info_rsc_dat_stride[31:0]),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .dma_read_ctrl_rsc_dat_size(dma_read_ctrl_rsc_dat_size),
      .dma_read_ctrl_rsc_dat_length(dma_read_ctrl_rsc_dat_length),
      .dma_read_ctrl_rsc_dat_index(dma_read_ctrl_rsc_dat_index),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_write_ctrl_rsc_dat_size(dma_write_ctrl_rsc_dat_size),
      .dma_write_ctrl_rsc_dat_length(dma_write_ctrl_rsc_dat_length),
      .dma_write_ctrl_rsc_dat_index(dma_write_ctrl_rsc_dat_index),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .acc_done_rsc_vld(acc_done_rsc_vld)
    );
  assign dma_read_ctrl_rsc_dat = {dma_read_ctrl_rsc_dat_size , dma_read_ctrl_rsc_dat_length
      , dma_read_ctrl_rsc_dat_index};
  assign dma_write_ctrl_rsc_dat = {dma_write_ctrl_rsc_dat_size , dma_write_ctrl_rsc_dat_length
      , dma_write_ctrl_rsc_dat_index};
endmodule



