
//------> ./conv2d_cxx_catapult_ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> ./conv2d_cxx_catapult_ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> ./conv2d_cxx_catapult_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2d_cxx_catapult_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> /tools/calypto/CATAPULT_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./conv2d_cxx_catapult.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   perenno@esp
//  Generated date: Mon Oct 31 22:08:01 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_9_14_32_10368_10368_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_9_14_32_10368_10368_32_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input clken_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_8_16_32_50176_50176_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_8_16_32_50176_50176_32_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [31:0] q;
  output [15:0] radr;
  output we;
  output [31:0] d;
  output [15:0] wadr;
  input clken_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [15:0] radr_d;
  input [15:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_7_14_32_10368_10368_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_7_14_32_10368_10368_32_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input clken_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_fsm (
  clk, rst, core_wen, fsm_output, BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input core_wen;
  output [3:0] fsm_output;
  reg [3:0] fsm_output;
  input BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_fsm_1
  parameter
    core_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    BATCH_LOOP_C_0 = 2'd2,
    main_C_1 = 2'd3;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 4'b0010;
        state_var_NS = BATCH_LOOP_C_0;
      end
      BATCH_LOOP_C_0 : begin
        fsm_output = 4'b0100;
        if ( BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = BATCH_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 4'b1000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 4'b0001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_staller (
  clk, rst, core_wen, core_wten, conf_info_rsci_wen_comp, dma_write_ctrl_rsci_wen_comp,
      dma_read_chnl_rsci_wen_comp, dma_write_chnl_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input conf_info_rsci_wen_comp;
  input dma_write_ctrl_rsci_wen_comp;
  input dma_read_chnl_rsci_wen_comp;
  input dma_write_chnl_rsci_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & dma_write_ctrl_rsci_wen_comp & dma_read_chnl_rsci_wen_comp
      & dma_write_chnl_rsci_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_dp
    (
  clk, rst, plm_out_data_rsci_q_d, plm_out_data_rsci_bawt, plm_out_data_rsci_q_d_mxwt,
      plm_out_data_rsci_biwt, plm_out_data_rsci_bdwt, plm_out_data_rsci_biwt_1, plm_out_data_rsci_bdwt_2
);
  input clk;
  input rst;
  input [31:0] plm_out_data_rsci_q_d;
  output plm_out_data_rsci_bawt;
  output [31:0] plm_out_data_rsci_q_d_mxwt;
  input plm_out_data_rsci_biwt;
  input plm_out_data_rsci_bdwt;
  input plm_out_data_rsci_biwt_1;
  input plm_out_data_rsci_bdwt_2;


  // Interconnect Declarations
  reg plm_out_data_rsci_bcwt;
  reg plm_out_data_rsci_bcwt_1;
  reg [31:0] plm_out_data_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_data_rsci_bawt = plm_out_data_rsci_biwt | plm_out_data_rsci_bcwt;
  assign plm_out_data_rsci_q_d_mxwt = MUX_v_32_2_2(plm_out_data_rsci_q_d, plm_out_data_rsci_q_d_bfwt,
      plm_out_data_rsci_bcwt_1);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_data_rsci_bcwt <= 1'b0;
      plm_out_data_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      plm_out_data_rsci_bcwt <= ~((~(plm_out_data_rsci_bcwt | plm_out_data_rsci_biwt))
          | plm_out_data_rsci_bdwt);
      plm_out_data_rsci_bcwt_1 <= ~((~(plm_out_data_rsci_bcwt_1 | plm_out_data_rsci_biwt_1))
          | plm_out_data_rsci_bdwt_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_data_rsci_q_d_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( plm_out_data_rsci_biwt_1 ) begin
      plm_out_data_rsci_q_d_bfwt <= plm_out_data_rsci_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_out_data_rsci_oswt_unreg, plm_out_data_rsci_iswt0, plm_out_data_rsci_oswt_unreg_1,
      plm_out_data_rsci_iswt0_1, plm_out_data_rsci_biwt, plm_out_data_rsci_bdwt,
      plm_out_data_rsci_biwt_1, plm_out_data_rsci_bdwt_2, plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct,
      plm_out_data_rsci_we_d_core_sct_pff, plm_out_data_rsci_iswt0_pff, plm_out_data_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input plm_out_data_rsci_oswt_unreg;
  input plm_out_data_rsci_iswt0;
  input plm_out_data_rsci_oswt_unreg_1;
  input plm_out_data_rsci_iswt0_1;
  output plm_out_data_rsci_biwt;
  output plm_out_data_rsci_bdwt;
  output plm_out_data_rsci_biwt_1;
  output plm_out_data_rsci_bdwt_2;
  output plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  output plm_out_data_rsci_we_d_core_sct_pff;
  input plm_out_data_rsci_iswt0_pff;
  input plm_out_data_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_data_rsci_bdwt = plm_out_data_rsci_oswt_unreg & core_wen;
  assign plm_out_data_rsci_biwt = (~ core_wten) & plm_out_data_rsci_iswt0;
  assign plm_out_data_rsci_bdwt_2 = plm_out_data_rsci_oswt_unreg_1 & core_wen;
  assign plm_out_data_rsci_biwt_1 = (~ core_wten) & plm_out_data_rsci_iswt0_1;
  assign plm_out_data_rsci_we_d_core_sct_pff = plm_out_data_rsci_iswt0_pff & core_wen;
  assign plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct = plm_out_data_rsci_iswt0_1_pff
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_dp
    (
  clk, rst, plm_f_data_rsci_q_d, plm_f_data_rsci_bawt, plm_f_data_rsci_q_d_mxwt,
      plm_f_data_rsci_biwt, plm_f_data_rsci_bdwt, plm_f_data_rsci_biwt_1, plm_f_data_rsci_bdwt_2
);
  input clk;
  input rst;
  input [31:0] plm_f_data_rsci_q_d;
  output plm_f_data_rsci_bawt;
  output [31:0] plm_f_data_rsci_q_d_mxwt;
  input plm_f_data_rsci_biwt;
  input plm_f_data_rsci_bdwt;
  input plm_f_data_rsci_biwt_1;
  input plm_f_data_rsci_bdwt_2;


  // Interconnect Declarations
  reg plm_f_data_rsci_bcwt;
  reg plm_f_data_rsci_bcwt_1;
  reg [31:0] plm_f_data_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_f_data_rsci_bawt = plm_f_data_rsci_biwt | plm_f_data_rsci_bcwt;
  assign plm_f_data_rsci_q_d_mxwt = MUX_v_32_2_2(plm_f_data_rsci_q_d, plm_f_data_rsci_q_d_bfwt,
      plm_f_data_rsci_bcwt_1);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_f_data_rsci_bcwt <= 1'b0;
      plm_f_data_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      plm_f_data_rsci_bcwt <= ~((~(plm_f_data_rsci_bcwt | plm_f_data_rsci_biwt))
          | plm_f_data_rsci_bdwt);
      plm_f_data_rsci_bcwt_1 <= ~((~(plm_f_data_rsci_bcwt_1 | plm_f_data_rsci_biwt_1))
          | plm_f_data_rsci_bdwt_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_f_data_rsci_q_d_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( plm_f_data_rsci_biwt_1 ) begin
      plm_f_data_rsci_q_d_bfwt <= plm_f_data_rsci_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_f_data_rsci_oswt_unreg, plm_f_data_rsci_iswt0, plm_f_data_rsci_oswt_unreg_1,
      plm_f_data_rsci_iswt0_1, plm_f_data_rsci_biwt, plm_f_data_rsci_bdwt, plm_f_data_rsci_biwt_1,
      plm_f_data_rsci_bdwt_2, plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct,
      plm_f_data_rsci_we_d_core_sct_pff, plm_f_data_rsci_iswt0_pff, plm_f_data_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input plm_f_data_rsci_oswt_unreg;
  input plm_f_data_rsci_iswt0;
  input plm_f_data_rsci_oswt_unreg_1;
  input plm_f_data_rsci_iswt0_1;
  output plm_f_data_rsci_biwt;
  output plm_f_data_rsci_bdwt;
  output plm_f_data_rsci_biwt_1;
  output plm_f_data_rsci_bdwt_2;
  output plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  output plm_f_data_rsci_we_d_core_sct_pff;
  input plm_f_data_rsci_iswt0_pff;
  input plm_f_data_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_f_data_rsci_bdwt = plm_f_data_rsci_oswt_unreg & core_wen;
  assign plm_f_data_rsci_biwt = (~ core_wten) & plm_f_data_rsci_iswt0;
  assign plm_f_data_rsci_bdwt_2 = plm_f_data_rsci_oswt_unreg_1 & core_wen;
  assign plm_f_data_rsci_biwt_1 = (~ core_wten) & plm_f_data_rsci_iswt0_1;
  assign plm_f_data_rsci_we_d_core_sct_pff = plm_f_data_rsci_iswt0_pff & core_wen;
  assign plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct = plm_f_data_rsci_iswt0_1_pff
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_dp
    (
  clk, rst, plm_in_data_rsci_q_d, plm_in_data_rsci_bawt, plm_in_data_rsci_q_d_mxwt,
      plm_in_data_rsci_biwt, plm_in_data_rsci_bdwt, plm_in_data_rsci_biwt_1, plm_in_data_rsci_bdwt_2
);
  input clk;
  input rst;
  input [31:0] plm_in_data_rsci_q_d;
  output plm_in_data_rsci_bawt;
  output [31:0] plm_in_data_rsci_q_d_mxwt;
  input plm_in_data_rsci_biwt;
  input plm_in_data_rsci_bdwt;
  input plm_in_data_rsci_biwt_1;
  input plm_in_data_rsci_bdwt_2;


  // Interconnect Declarations
  reg plm_in_data_rsci_bcwt;
  reg plm_in_data_rsci_bcwt_1;
  reg [31:0] plm_in_data_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_data_rsci_bawt = plm_in_data_rsci_biwt | plm_in_data_rsci_bcwt;
  assign plm_in_data_rsci_q_d_mxwt = MUX_v_32_2_2(plm_in_data_rsci_q_d, plm_in_data_rsci_q_d_bfwt,
      plm_in_data_rsci_bcwt_1);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_data_rsci_bcwt <= 1'b0;
      plm_in_data_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      plm_in_data_rsci_bcwt <= ~((~(plm_in_data_rsci_bcwt | plm_in_data_rsci_biwt))
          | plm_in_data_rsci_bdwt);
      plm_in_data_rsci_bcwt_1 <= ~((~(plm_in_data_rsci_bcwt_1 | plm_in_data_rsci_biwt_1))
          | plm_in_data_rsci_bdwt_2);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_data_rsci_q_d_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( plm_in_data_rsci_biwt_1 ) begin
      plm_in_data_rsci_q_d_bfwt <= plm_in_data_rsci_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_in_data_rsci_oswt_unreg, plm_in_data_rsci_iswt0, plm_in_data_rsci_oswt_unreg_1,
      plm_in_data_rsci_iswt0_1, plm_in_data_rsci_biwt, plm_in_data_rsci_bdwt, plm_in_data_rsci_biwt_1,
      plm_in_data_rsci_bdwt_2, plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct,
      plm_in_data_rsci_we_d_core_sct_pff, plm_in_data_rsci_iswt0_pff, plm_in_data_rsci_iswt0_1_pff
);
  input core_wen;
  input core_wten;
  input plm_in_data_rsci_oswt_unreg;
  input plm_in_data_rsci_iswt0;
  input plm_in_data_rsci_oswt_unreg_1;
  input plm_in_data_rsci_iswt0_1;
  output plm_in_data_rsci_biwt;
  output plm_in_data_rsci_bdwt;
  output plm_in_data_rsci_biwt_1;
  output plm_in_data_rsci_bdwt_2;
  output plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  output plm_in_data_rsci_we_d_core_sct_pff;
  input plm_in_data_rsci_iswt0_pff;
  input plm_in_data_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_data_rsci_bdwt = plm_in_data_rsci_oswt_unreg & core_wen;
  assign plm_in_data_rsci_biwt = (~ core_wten) & plm_in_data_rsci_iswt0;
  assign plm_in_data_rsci_bdwt_2 = plm_in_data_rsci_oswt_unreg_1 & core_wen;
  assign plm_in_data_rsci_biwt_1 = (~ core_wten) & plm_in_data_rsci_iswt0_1;
  assign plm_in_data_rsci_we_d_core_sct_pff = plm_in_data_rsci_iswt0_pff & core_wen;
  assign plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct = plm_in_data_rsci_iswt0_1_pff
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_acc_done_rsci_acc_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_acc_done_rsci_acc_done_wait_ctrl
    (
  core_wten, acc_done_rsci_iswt0, acc_done_rsci_ivld_core_sct
);
  input core_wten;
  input acc_done_rsci_iswt0;
  output acc_done_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign acc_done_rsci_ivld_core_sct = acc_done_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
    (
  clk, rst, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_bawt, dma_write_chnl_rsci_wen_comp,
      dma_write_chnl_rsci_biwt, dma_write_chnl_rsci_bdwt, dma_write_chnl_rsci_bcwt
);
  input clk;
  input rst;
  input dma_write_chnl_rsci_oswt_unreg;
  output dma_write_chnl_rsci_bawt;
  output dma_write_chnl_rsci_wen_comp;
  input dma_write_chnl_rsci_biwt;
  input dma_write_chnl_rsci_bdwt;
  output dma_write_chnl_rsci_bcwt;
  reg dma_write_chnl_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_rsci_bawt = dma_write_chnl_rsci_biwt | dma_write_chnl_rsci_bcwt;
  assign dma_write_chnl_rsci_wen_comp = (~ dma_write_chnl_rsci_oswt_unreg) | dma_write_chnl_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_write_chnl_rsci_bcwt <= ~((~(dma_write_chnl_rsci_bcwt | dma_write_chnl_rsci_biwt))
          | dma_write_chnl_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
    (
  core_wen, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_iswt0, dma_write_chnl_rsci_irdy,
      dma_write_chnl_rsci_biwt, dma_write_chnl_rsci_bdwt, dma_write_chnl_rsci_bcwt,
      dma_write_chnl_rsci_ivld_core_sct
);
  input core_wen;
  input dma_write_chnl_rsci_oswt_unreg;
  input dma_write_chnl_rsci_iswt0;
  input dma_write_chnl_rsci_irdy;
  output dma_write_chnl_rsci_biwt;
  output dma_write_chnl_rsci_bdwt;
  input dma_write_chnl_rsci_bcwt;
  output dma_write_chnl_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire dma_write_chnl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_rsci_bdwt = dma_write_chnl_rsci_oswt_unreg & core_wen;
  assign dma_write_chnl_rsci_biwt = dma_write_chnl_rsci_ogwt & dma_write_chnl_rsci_irdy;
  assign dma_write_chnl_rsci_ogwt = dma_write_chnl_rsci_iswt0 & (~ dma_write_chnl_rsci_bcwt);
  assign dma_write_chnl_rsci_ivld_core_sct = dma_write_chnl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
    (
  clk, rst, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_bawt, dma_read_chnl_rsci_wen_comp,
      dma_read_chnl_rsci_idat_mxwt, dma_read_chnl_rsci_biwt, dma_read_chnl_rsci_bdwt,
      dma_read_chnl_rsci_bcwt, dma_read_chnl_rsci_idat
);
  input clk;
  input rst;
  input dma_read_chnl_rsci_oswt_unreg;
  output dma_read_chnl_rsci_bawt;
  output dma_read_chnl_rsci_wen_comp;
  output [31:0] dma_read_chnl_rsci_idat_mxwt;
  input dma_read_chnl_rsci_biwt;
  input dma_read_chnl_rsci_bdwt;
  output dma_read_chnl_rsci_bcwt;
  reg dma_read_chnl_rsci_bcwt;
  input [63:0] dma_read_chnl_rsci_idat;


  // Interconnect Declarations
  reg [31:0] dma_read_chnl_rsci_idat_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_rsci_bawt = dma_read_chnl_rsci_biwt | dma_read_chnl_rsci_bcwt;
  assign dma_read_chnl_rsci_wen_comp = (~ dma_read_chnl_rsci_oswt_unreg) | dma_read_chnl_rsci_bawt;
  assign dma_read_chnl_rsci_idat_mxwt = MUX_v_32_2_2((dma_read_chnl_rsci_idat[31:0]),
      dma_read_chnl_rsci_idat_bfwt_31_0, dma_read_chnl_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_read_chnl_rsci_bcwt <= ~((~(dma_read_chnl_rsci_bcwt | dma_read_chnl_rsci_biwt))
          | dma_read_chnl_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_rsci_idat_bfwt_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( dma_read_chnl_rsci_biwt ) begin
      dma_read_chnl_rsci_idat_bfwt_31_0 <= dma_read_chnl_rsci_idat[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
    (
  core_wen, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_iswt0, dma_read_chnl_rsci_biwt,
      dma_read_chnl_rsci_bdwt, dma_read_chnl_rsci_bcwt, dma_read_chnl_rsci_irdy_core_sct,
      dma_read_chnl_rsci_ivld
);
  input core_wen;
  input dma_read_chnl_rsci_oswt_unreg;
  input dma_read_chnl_rsci_iswt0;
  output dma_read_chnl_rsci_biwt;
  output dma_read_chnl_rsci_bdwt;
  input dma_read_chnl_rsci_bcwt;
  output dma_read_chnl_rsci_irdy_core_sct;
  input dma_read_chnl_rsci_ivld;


  // Interconnect Declarations
  wire dma_read_chnl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_rsci_bdwt = dma_read_chnl_rsci_oswt_unreg & core_wen;
  assign dma_read_chnl_rsci_biwt = dma_read_chnl_rsci_ogwt & dma_read_chnl_rsci_ivld;
  assign dma_read_chnl_rsci_ogwt = dma_read_chnl_rsci_iswt0 & (~ dma_read_chnl_rsci_bcwt);
  assign dma_read_chnl_rsci_irdy_core_sct = dma_read_chnl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
    (
  clk, rst, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_bawt, dma_write_ctrl_rsci_wen_comp,
      dma_write_ctrl_rsci_biwt, dma_write_ctrl_rsci_bdwt, dma_write_ctrl_rsci_bcwt
);
  input clk;
  input rst;
  input dma_write_ctrl_rsci_oswt_unreg;
  output dma_write_ctrl_rsci_bawt;
  output dma_write_ctrl_rsci_wen_comp;
  input dma_write_ctrl_rsci_biwt;
  input dma_write_ctrl_rsci_bdwt;
  output dma_write_ctrl_rsci_bcwt;
  reg dma_write_ctrl_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_rsci_bawt = dma_write_ctrl_rsci_biwt | dma_write_ctrl_rsci_bcwt;
  assign dma_write_ctrl_rsci_wen_comp = (~ dma_write_ctrl_rsci_oswt_unreg) | dma_write_ctrl_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_rsci_bcwt <= ~((~(dma_write_ctrl_rsci_bcwt | dma_write_ctrl_rsci_biwt))
          | dma_write_ctrl_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
    (
  core_wen, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_iswt0, dma_write_ctrl_rsci_irdy,
      dma_write_ctrl_rsci_biwt, dma_write_ctrl_rsci_bdwt, dma_write_ctrl_rsci_bcwt,
      dma_write_ctrl_rsci_ivld_core_sct
);
  input core_wen;
  input dma_write_ctrl_rsci_oswt_unreg;
  input dma_write_ctrl_rsci_iswt0;
  input dma_write_ctrl_rsci_irdy;
  output dma_write_ctrl_rsci_biwt;
  output dma_write_ctrl_rsci_bdwt;
  input dma_write_ctrl_rsci_bcwt;
  output dma_write_ctrl_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire dma_write_ctrl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_rsci_bdwt = dma_write_ctrl_rsci_oswt_unreg & core_wen;
  assign dma_write_ctrl_rsci_biwt = dma_write_ctrl_rsci_ogwt & dma_write_ctrl_rsci_irdy;
  assign dma_write_ctrl_rsci_ogwt = dma_write_ctrl_rsci_iswt0 & (~ dma_write_ctrl_rsci_bcwt);
  assign dma_write_ctrl_rsci_ivld_core_sct = dma_write_ctrl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
    (
  clk, rst, dma_read_ctrl_rsci_bawt, dma_read_ctrl_rsci_irdy_mxwt, dma_read_ctrl_rsci_irdy,
      dma_read_ctrl_rsci_biwt, dma_read_ctrl_rsci_bdwt
);
  input clk;
  input rst;
  output dma_read_ctrl_rsci_bawt;
  output dma_read_ctrl_rsci_irdy_mxwt;
  input dma_read_ctrl_rsci_irdy;
  input dma_read_ctrl_rsci_biwt;
  input dma_read_ctrl_rsci_bdwt;


  // Interconnect Declarations
  reg dma_read_ctrl_rsci_bcwt;
  reg dma_read_ctrl_rsci_irdy_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_rsci_bawt = dma_read_ctrl_rsci_biwt | dma_read_ctrl_rsci_bcwt;
  assign dma_read_ctrl_rsci_irdy_mxwt = MUX_s_1_2_2(dma_read_ctrl_rsci_irdy, dma_read_ctrl_rsci_irdy_bfwt,
      dma_read_ctrl_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_rsci_bcwt <= ~((~(dma_read_ctrl_rsci_bcwt | dma_read_ctrl_rsci_biwt))
          | dma_read_ctrl_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_irdy_bfwt <= 1'b0;
    end
    else if ( dma_read_ctrl_rsci_biwt ) begin
      dma_read_ctrl_rsci_irdy_bfwt <= dma_read_ctrl_rsci_irdy;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
    (
  core_wen, core_wten, dma_read_ctrl_rsci_oswt_unreg, dma_read_ctrl_rsci_iswt0, dma_read_ctrl_rsci_biwt,
      dma_read_ctrl_rsci_bdwt
);
  input core_wen;
  input core_wten;
  input dma_read_ctrl_rsci_oswt_unreg;
  input dma_read_ctrl_rsci_iswt0;
  output dma_read_ctrl_rsci_biwt;
  output dma_read_ctrl_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_rsci_bdwt = dma_read_ctrl_rsci_oswt_unreg & core_wen;
  assign dma_read_ctrl_rsci_biwt = (~ core_wten) & dma_read_ctrl_rsci_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_dp
    (
  clk, rst, conf_info_rsci_oswt, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt,
      conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt;
  output conf_info_rsci_wen_comp;
  output [231:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  reg [231:0] conf_info_rsci_idat_bfwt_231_0;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt) | conf_info_rsci_biwt
      | conf_info_rsci_bcwt;
  assign conf_info_rsci_idat_mxwt = MUX_v_232_2_2((conf_info_rsci_idat[231:0]), conf_info_rsci_idat_bfwt_231_0,
      conf_info_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt_231_0 <= conf_info_rsci_idat[231:0];
    end
  end

  function automatic [231:0] MUX_v_232_2_2;
    input [231:0] input_0;
    input [231:0] input_1;
    input [0:0] sel;
    reg [231:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_232_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_oswt & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1 (
  clk, rst, plm_out_data_rsci_q_d, plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, plm_out_data_rsci_oswt_unreg, plm_out_data_rsci_bawt,
      plm_out_data_rsci_iswt0, plm_out_data_rsci_oswt_unreg_1, plm_out_data_rsci_iswt0_1,
      plm_out_data_rsci_q_d_mxwt, plm_out_data_rsci_we_d_pff, plm_out_data_rsci_iswt0_pff,
      plm_out_data_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  input [31:0] plm_out_data_rsci_q_d;
  output plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input plm_out_data_rsci_oswt_unreg;
  output plm_out_data_rsci_bawt;
  input plm_out_data_rsci_iswt0;
  input plm_out_data_rsci_oswt_unreg_1;
  input plm_out_data_rsci_iswt0_1;
  output [31:0] plm_out_data_rsci_q_d_mxwt;
  output plm_out_data_rsci_we_d_pff;
  input plm_out_data_rsci_iswt0_pff;
  input plm_out_data_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire plm_out_data_rsci_biwt;
  wire plm_out_data_rsci_bdwt;
  wire plm_out_data_rsci_biwt_1;
  wire plm_out_data_rsci_bdwt_2;
  wire plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  wire plm_out_data_rsci_we_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_ctrl
      conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_out_data_rsci_oswt_unreg(plm_out_data_rsci_oswt_unreg),
      .plm_out_data_rsci_iswt0(plm_out_data_rsci_iswt0),
      .plm_out_data_rsci_oswt_unreg_1(plm_out_data_rsci_oswt_unreg_1),
      .plm_out_data_rsci_iswt0_1(plm_out_data_rsci_iswt0_1),
      .plm_out_data_rsci_biwt(plm_out_data_rsci_biwt),
      .plm_out_data_rsci_bdwt(plm_out_data_rsci_bdwt),
      .plm_out_data_rsci_biwt_1(plm_out_data_rsci_biwt_1),
      .plm_out_data_rsci_bdwt_2(plm_out_data_rsci_bdwt_2),
      .plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct(plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct),
      .plm_out_data_rsci_we_d_core_sct_pff(plm_out_data_rsci_we_d_core_sct_iff),
      .plm_out_data_rsci_iswt0_pff(plm_out_data_rsci_iswt0_pff),
      .plm_out_data_rsci_iswt0_1_pff(plm_out_data_rsci_iswt0_1_pff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_dp
      conv2d_cxx_catapult_core_plm_out_data_rsci_1_plm_out_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_data_rsci_q_d(plm_out_data_rsci_q_d),
      .plm_out_data_rsci_bawt(plm_out_data_rsci_bawt),
      .plm_out_data_rsci_q_d_mxwt(plm_out_data_rsci_q_d_mxwt),
      .plm_out_data_rsci_biwt(plm_out_data_rsci_biwt),
      .plm_out_data_rsci_bdwt(plm_out_data_rsci_bdwt),
      .plm_out_data_rsci_biwt_1(plm_out_data_rsci_biwt_1),
      .plm_out_data_rsci_bdwt_2(plm_out_data_rsci_bdwt_2)
    );
  assign plm_out_data_rsci_we_d_pff = plm_out_data_rsci_we_d_core_sct_iff;
  assign plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1 (
  clk, rst, plm_f_data_rsci_q_d, plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, plm_f_data_rsci_oswt_unreg, plm_f_data_rsci_bawt, plm_f_data_rsci_iswt0,
      plm_f_data_rsci_oswt_unreg_1, plm_f_data_rsci_iswt0_1, plm_f_data_rsci_q_d_mxwt,
      plm_f_data_rsci_we_d_pff, plm_f_data_rsci_iswt0_pff, plm_f_data_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  input [31:0] plm_f_data_rsci_q_d;
  output plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input plm_f_data_rsci_oswt_unreg;
  output plm_f_data_rsci_bawt;
  input plm_f_data_rsci_iswt0;
  input plm_f_data_rsci_oswt_unreg_1;
  input plm_f_data_rsci_iswt0_1;
  output [31:0] plm_f_data_rsci_q_d_mxwt;
  output plm_f_data_rsci_we_d_pff;
  input plm_f_data_rsci_iswt0_pff;
  input plm_f_data_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire plm_f_data_rsci_biwt;
  wire plm_f_data_rsci_bdwt;
  wire plm_f_data_rsci_biwt_1;
  wire plm_f_data_rsci_bdwt_2;
  wire plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  wire plm_f_data_rsci_we_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_ctrl
      conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_f_data_rsci_oswt_unreg(plm_f_data_rsci_oswt_unreg),
      .plm_f_data_rsci_iswt0(plm_f_data_rsci_iswt0),
      .plm_f_data_rsci_oswt_unreg_1(plm_f_data_rsci_oswt_unreg_1),
      .plm_f_data_rsci_iswt0_1(plm_f_data_rsci_iswt0_1),
      .plm_f_data_rsci_biwt(plm_f_data_rsci_biwt),
      .plm_f_data_rsci_bdwt(plm_f_data_rsci_bdwt),
      .plm_f_data_rsci_biwt_1(plm_f_data_rsci_biwt_1),
      .plm_f_data_rsci_bdwt_2(plm_f_data_rsci_bdwt_2),
      .plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct(plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct),
      .plm_f_data_rsci_we_d_core_sct_pff(plm_f_data_rsci_we_d_core_sct_iff),
      .plm_f_data_rsci_iswt0_pff(plm_f_data_rsci_iswt0_pff),
      .plm_f_data_rsci_iswt0_1_pff(plm_f_data_rsci_iswt0_1_pff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_dp
      conv2d_cxx_catapult_core_plm_f_data_rsci_1_plm_f_data_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_f_data_rsci_q_d(plm_f_data_rsci_q_d),
      .plm_f_data_rsci_bawt(plm_f_data_rsci_bawt),
      .plm_f_data_rsci_q_d_mxwt(plm_f_data_rsci_q_d_mxwt),
      .plm_f_data_rsci_biwt(plm_f_data_rsci_biwt),
      .plm_f_data_rsci_bdwt(plm_f_data_rsci_bdwt),
      .plm_f_data_rsci_biwt_1(plm_f_data_rsci_biwt_1),
      .plm_f_data_rsci_bdwt_2(plm_f_data_rsci_bdwt_2)
    );
  assign plm_f_data_rsci_we_d_pff = plm_f_data_rsci_we_d_core_sct_iff;
  assign plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1 (
  clk, rst, plm_in_data_rsci_q_d, plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, plm_in_data_rsci_oswt_unreg, plm_in_data_rsci_bawt, plm_in_data_rsci_iswt0,
      plm_in_data_rsci_oswt_unreg_1, plm_in_data_rsci_iswt0_1, plm_in_data_rsci_q_d_mxwt,
      plm_in_data_rsci_we_d_pff, plm_in_data_rsci_iswt0_pff, plm_in_data_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  input [31:0] plm_in_data_rsci_q_d;
  output plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input plm_in_data_rsci_oswt_unreg;
  output plm_in_data_rsci_bawt;
  input plm_in_data_rsci_iswt0;
  input plm_in_data_rsci_oswt_unreg_1;
  input plm_in_data_rsci_iswt0_1;
  output [31:0] plm_in_data_rsci_q_d_mxwt;
  output plm_in_data_rsci_we_d_pff;
  input plm_in_data_rsci_iswt0_pff;
  input plm_in_data_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire plm_in_data_rsci_biwt;
  wire plm_in_data_rsci_bdwt;
  wire plm_in_data_rsci_biwt_1;
  wire plm_in_data_rsci_bdwt_2;
  wire plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  wire plm_in_data_rsci_we_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_ctrl
      conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_in_data_rsci_oswt_unreg(plm_in_data_rsci_oswt_unreg),
      .plm_in_data_rsci_iswt0(plm_in_data_rsci_iswt0),
      .plm_in_data_rsci_oswt_unreg_1(plm_in_data_rsci_oswt_unreg_1),
      .plm_in_data_rsci_iswt0_1(plm_in_data_rsci_iswt0_1),
      .plm_in_data_rsci_biwt(plm_in_data_rsci_biwt),
      .plm_in_data_rsci_bdwt(plm_in_data_rsci_bdwt),
      .plm_in_data_rsci_biwt_1(plm_in_data_rsci_biwt_1),
      .plm_in_data_rsci_bdwt_2(plm_in_data_rsci_bdwt_2),
      .plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct(plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct),
      .plm_in_data_rsci_we_d_core_sct_pff(plm_in_data_rsci_we_d_core_sct_iff),
      .plm_in_data_rsci_iswt0_pff(plm_in_data_rsci_iswt0_pff),
      .plm_in_data_rsci_iswt0_1_pff(plm_in_data_rsci_iswt0_1_pff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_dp
      conv2d_cxx_catapult_core_plm_in_data_rsci_1_plm_in_data_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_in_data_rsci_q_d(plm_in_data_rsci_q_d),
      .plm_in_data_rsci_bawt(plm_in_data_rsci_bawt),
      .plm_in_data_rsci_q_d_mxwt(plm_in_data_rsci_q_d_mxwt),
      .plm_in_data_rsci_biwt(plm_in_data_rsci_biwt),
      .plm_in_data_rsci_bdwt(plm_in_data_rsci_bdwt),
      .plm_in_data_rsci_biwt_1(plm_in_data_rsci_biwt_1),
      .plm_in_data_rsci_bdwt_2(plm_in_data_rsci_bdwt_2)
    );
  assign plm_in_data_rsci_we_d_pff = plm_in_data_rsci_we_d_core_sct_iff;
  assign plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_acc_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_acc_done_rsci (
  acc_done_rsc_vld, core_wten, acc_done_rsci_iswt0
);
  output acc_done_rsc_vld;
  input core_wten;
  input acc_done_rsci_iswt0;


  // Interconnect Declarations
  wire acc_done_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_out_vld_v1 #(.rscid(32'sd6)) acc_done_rsci
      (
      .vld(acc_done_rsc_vld),
      .ivld(acc_done_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_acc_done_rsci_acc_done_wait_ctrl
      conv2d_cxx_catapult_core_acc_done_rsci_acc_done_wait_ctrl_inst (
      .core_wten(core_wten),
      .acc_done_rsci_iswt0(acc_done_rsci_iswt0),
      .acc_done_rsci_ivld_core_sct(acc_done_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci (
  clk, rst, dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy,
      core_wen, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_bawt, dma_write_chnl_rsci_iswt0,
      dma_write_chnl_rsci_wen_comp, dma_write_chnl_rsci_idat
);
  input clk;
  input rst;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  input core_wen;
  input dma_write_chnl_rsci_oswt_unreg;
  output dma_write_chnl_rsci_bawt;
  input dma_write_chnl_rsci_iswt0;
  output dma_write_chnl_rsci_wen_comp;
  input [63:0] dma_write_chnl_rsci_idat;


  // Interconnect Declarations
  wire dma_write_chnl_rsci_irdy;
  wire dma_write_chnl_rsci_biwt;
  wire dma_write_chnl_rsci_bdwt;
  wire dma_write_chnl_rsci_bcwt;
  wire dma_write_chnl_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_dma_write_chnl_rsci_idat;
  assign nl_dma_write_chnl_rsci_idat = {32'b11011110101011011011111011101111 , (dma_write_chnl_rsci_idat[31:0])};
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd5),
  .width(32'sd64)) dma_write_chnl_rsci (
      .irdy(dma_write_chnl_rsci_irdy),
      .ivld(dma_write_chnl_rsci_ivld_core_sct),
      .idat(nl_dma_write_chnl_rsci_idat[63:0]),
      .rdy(dma_write_chnl_rsc_rdy),
      .vld(dma_write_chnl_rsc_vld),
      .dat(dma_write_chnl_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
      conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .dma_write_chnl_rsci_oswt_unreg(dma_write_chnl_rsci_oswt_unreg),
      .dma_write_chnl_rsci_iswt0(dma_write_chnl_rsci_iswt0),
      .dma_write_chnl_rsci_irdy(dma_write_chnl_rsci_irdy),
      .dma_write_chnl_rsci_biwt(dma_write_chnl_rsci_biwt),
      .dma_write_chnl_rsci_bdwt(dma_write_chnl_rsci_bdwt),
      .dma_write_chnl_rsci_bcwt(dma_write_chnl_rsci_bcwt),
      .dma_write_chnl_rsci_ivld_core_sct(dma_write_chnl_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
      conv2d_cxx_catapult_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_rsci_oswt_unreg(dma_write_chnl_rsci_oswt_unreg),
      .dma_write_chnl_rsci_bawt(dma_write_chnl_rsci_bawt),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .dma_write_chnl_rsci_biwt(dma_write_chnl_rsci_biwt),
      .dma_write_chnl_rsci_bdwt(dma_write_chnl_rsci_bdwt),
      .dma_write_chnl_rsci_bcwt(dma_write_chnl_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci (
  clk, rst, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy,
      core_wen, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_bawt, dma_read_chnl_rsci_iswt0,
      dma_read_chnl_rsci_wen_comp, dma_read_chnl_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  input core_wen;
  input dma_read_chnl_rsci_oswt_unreg;
  output dma_read_chnl_rsci_bawt;
  input dma_read_chnl_rsci_iswt0;
  output dma_read_chnl_rsci_wen_comp;
  output [31:0] dma_read_chnl_rsci_idat_mxwt;


  // Interconnect Declarations
  wire dma_read_chnl_rsci_biwt;
  wire dma_read_chnl_rsci_bdwt;
  wire dma_read_chnl_rsci_bcwt;
  wire dma_read_chnl_rsci_irdy_core_sct;
  wire dma_read_chnl_rsci_ivld;
  wire [63:0] dma_read_chnl_rsci_idat;
  wire [31:0] dma_read_chnl_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd4),
  .width(32'sd64)) dma_read_chnl_rsci (
      .rdy(dma_read_chnl_rsc_rdy),
      .vld(dma_read_chnl_rsc_vld),
      .dat(dma_read_chnl_rsc_dat),
      .irdy(dma_read_chnl_rsci_irdy_core_sct),
      .ivld(dma_read_chnl_rsci_ivld),
      .idat(dma_read_chnl_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
      conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl_inst (
      .core_wen(core_wen),
      .dma_read_chnl_rsci_oswt_unreg(dma_read_chnl_rsci_oswt_unreg),
      .dma_read_chnl_rsci_iswt0(dma_read_chnl_rsci_iswt0),
      .dma_read_chnl_rsci_biwt(dma_read_chnl_rsci_biwt),
      .dma_read_chnl_rsci_bdwt(dma_read_chnl_rsci_bdwt),
      .dma_read_chnl_rsci_bcwt(dma_read_chnl_rsci_bcwt),
      .dma_read_chnl_rsci_irdy_core_sct(dma_read_chnl_rsci_irdy_core_sct),
      .dma_read_chnl_rsci_ivld(dma_read_chnl_rsci_ivld)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
      conv2d_cxx_catapult_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_rsci_oswt_unreg(dma_read_chnl_rsci_oswt_unreg),
      .dma_read_chnl_rsci_bawt(dma_read_chnl_rsci_bawt),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .dma_read_chnl_rsci_idat_mxwt(dma_read_chnl_rsci_idat_mxwt_pconst),
      .dma_read_chnl_rsci_biwt(dma_read_chnl_rsci_biwt),
      .dma_read_chnl_rsci_bdwt(dma_read_chnl_rsci_bdwt),
      .dma_read_chnl_rsci_bcwt(dma_read_chnl_rsci_bcwt),
      .dma_read_chnl_rsci_idat(dma_read_chnl_rsci_idat)
    );
  assign dma_read_chnl_rsci_idat_mxwt = dma_read_chnl_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci (
  clk, rst, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy,
      core_wen, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_bawt, dma_write_ctrl_rsci_iswt0,
      dma_write_ctrl_rsci_wen_comp, dma_write_ctrl_rsci_idat
);
  input clk;
  input rst;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input core_wen;
  input dma_write_ctrl_rsci_oswt_unreg;
  output dma_write_ctrl_rsci_bawt;
  input dma_write_ctrl_rsci_iswt0;
  output dma_write_ctrl_rsci_wen_comp;
  input [66:0] dma_write_ctrl_rsci_idat;


  // Interconnect Declarations
  wire dma_write_ctrl_rsci_irdy;
  wire dma_write_ctrl_rsci_biwt;
  wire dma_write_ctrl_rsci_bdwt;
  wire dma_write_ctrl_rsci_bcwt;
  wire dma_write_ctrl_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [66:0] nl_dma_write_ctrl_rsci_idat;
  assign nl_dma_write_ctrl_rsci_idat = {19'b0110000000000000000 , (dma_write_ctrl_rsci_idat[47:32])
      , 16'b0000000000000000 , (dma_write_ctrl_rsci_idat[15:0])};
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd67)) dma_write_ctrl_rsci (
      .irdy(dma_write_ctrl_rsci_irdy),
      .ivld(dma_write_ctrl_rsci_ivld_core_sct),
      .idat(nl_dma_write_ctrl_rsci_idat[66:0]),
      .rdy(dma_write_ctrl_rsc_rdy),
      .vld(dma_write_ctrl_rsc_vld),
      .dat(dma_write_ctrl_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
      conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .dma_write_ctrl_rsci_oswt_unreg(dma_write_ctrl_rsci_oswt_unreg),
      .dma_write_ctrl_rsci_iswt0(dma_write_ctrl_rsci_iswt0),
      .dma_write_ctrl_rsci_irdy(dma_write_ctrl_rsci_irdy),
      .dma_write_ctrl_rsci_biwt(dma_write_ctrl_rsci_biwt),
      .dma_write_ctrl_rsci_bdwt(dma_write_ctrl_rsci_bdwt),
      .dma_write_ctrl_rsci_bcwt(dma_write_ctrl_rsci_bcwt),
      .dma_write_ctrl_rsci_ivld_core_sct(dma_write_ctrl_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
      conv2d_cxx_catapult_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_rsci_oswt_unreg(dma_write_ctrl_rsci_oswt_unreg),
      .dma_write_ctrl_rsci_bawt(dma_write_ctrl_rsci_bawt),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_ctrl_rsci_biwt(dma_write_ctrl_rsci_biwt),
      .dma_write_ctrl_rsci_bdwt(dma_write_ctrl_rsci_bdwt),
      .dma_write_ctrl_rsci_bcwt(dma_write_ctrl_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci (
  clk, rst, dma_read_ctrl_rsc_dat, dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy,
      core_wen, core_wten, dma_read_ctrl_rsci_oswt_unreg, dma_read_ctrl_rsci_bawt,
      dma_read_ctrl_rsci_iswt0, dma_read_ctrl_rsci_irdy_mxwt, dma_read_ctrl_rsci_idat
);
  input clk;
  input rst;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  input core_wen;
  input core_wten;
  input dma_read_ctrl_rsci_oswt_unreg;
  output dma_read_ctrl_rsci_bawt;
  input dma_read_ctrl_rsci_iswt0;
  output dma_read_ctrl_rsci_irdy_mxwt;
  input [66:0] dma_read_ctrl_rsci_idat;


  // Interconnect Declarations
  wire dma_read_ctrl_rsci_irdy;
  wire dma_read_ctrl_rsci_biwt;
  wire dma_read_ctrl_rsci_bdwt;


  // Interconnect Declarations for Component Instantiations 
  wire [66:0] nl_dma_read_ctrl_rsci_idat;
  assign nl_dma_read_ctrl_rsci_idat = {19'b0110000000000000000 , (dma_read_ctrl_rsci_idat[47:32])
      , 16'b0000000000000000 , (dma_read_ctrl_rsci_idat[15:0])};
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd67)) dma_read_ctrl_rsci (
      .irdy(dma_read_ctrl_rsci_irdy),
      .ivld(dma_read_ctrl_rsci_biwt),
      .idat(nl_dma_read_ctrl_rsci_idat[66:0]),
      .rdy(dma_read_ctrl_rsc_rdy),
      .vld(dma_read_ctrl_rsc_vld),
      .dat(dma_read_ctrl_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
      conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dma_read_ctrl_rsci_oswt_unreg(dma_read_ctrl_rsci_oswt_unreg),
      .dma_read_ctrl_rsci_iswt0(dma_read_ctrl_rsci_iswt0),
      .dma_read_ctrl_rsci_biwt(dma_read_ctrl_rsci_biwt),
      .dma_read_ctrl_rsci_bdwt(dma_read_ctrl_rsci_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
      conv2d_cxx_catapult_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_rsci_bawt(dma_read_ctrl_rsci_bawt),
      .dma_read_ctrl_rsci_irdy_mxwt(dma_read_ctrl_rsci_irdy_mxwt),
      .dma_read_ctrl_rsci_irdy(dma_read_ctrl_rsci_irdy),
      .dma_read_ctrl_rsci_biwt(dma_read_ctrl_rsci_biwt),
      .dma_read_ctrl_rsci_bdwt(dma_read_ctrl_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt,
      conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt;
  output conf_info_rsci_wen_comp;
  output [231:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;
  wire [231:0] conf_info_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_ctrl
      conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_ctrl_inst (
      .core_wen(core_wen),
      .conf_info_rsci_oswt(conf_info_rsci_oswt),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_dp
      conv2d_cxx_catapult_core_conf_info_rsci_conf_info_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt(conf_info_rsci_oswt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt_pconst),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
  assign conf_info_rsci_idat_mxwt = conf_info_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, dma_read_ctrl_rsc_dat,
      dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld,
      dma_write_ctrl_rsc_rdy, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy,
      dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, acc_done_rsc_vld,
      plm_in_data_rsci_d_d, plm_in_data_rsci_q_d, plm_in_data_rsci_radr_d, plm_in_data_rsci_wadr_d,
      plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d, plm_f_data_rsci_d_d, plm_f_data_rsci_q_d,
      plm_f_data_rsci_radr_d, plm_f_data_rsci_wadr_d, plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      plm_out_data_rsci_d_d, plm_out_data_rsci_q_d, plm_out_data_rsci_radr_d, plm_out_data_rsci_wadr_d,
      plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d, plm_in_data_rsci_we_d_pff,
      plm_f_data_rsci_we_d_pff, plm_out_data_rsci_we_d_pff
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  output acc_done_rsc_vld;
  output [31:0] plm_in_data_rsci_d_d;
  input [31:0] plm_in_data_rsci_q_d;
  output [13:0] plm_in_data_rsci_radr_d;
  output [13:0] plm_in_data_rsci_wadr_d;
  output plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output [31:0] plm_f_data_rsci_d_d;
  input [31:0] plm_f_data_rsci_q_d;
  output [15:0] plm_f_data_rsci_radr_d;
  output [15:0] plm_f_data_rsci_wadr_d;
  output plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output [31:0] plm_out_data_rsci_d_d;
  input [31:0] plm_out_data_rsci_q_d;
  output [13:0] plm_out_data_rsci_radr_d;
  output [13:0] plm_out_data_rsci_wadr_d;
  output plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output plm_in_data_rsci_we_d_pff;
  output plm_f_data_rsci_we_d_pff;
  output plm_out_data_rsci_we_d_pff;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire conf_info_rsci_wen_comp;
  wire [231:0] conf_info_rsci_idat_mxwt;
  wire dma_read_ctrl_rsci_bawt;
  wire dma_read_ctrl_rsci_irdy_mxwt;
  wire dma_write_ctrl_rsci_bawt;
  wire dma_write_ctrl_rsci_wen_comp;
  wire dma_read_chnl_rsci_bawt;
  wire dma_read_chnl_rsci_wen_comp;
  wire [31:0] dma_read_chnl_rsci_idat_mxwt;
  wire dma_write_chnl_rsci_bawt;
  wire dma_write_chnl_rsci_wen_comp;
  wire plm_in_data_rsci_bawt;
  wire [31:0] plm_in_data_rsci_q_d_mxwt;
  wire plm_f_data_rsci_bawt;
  wire [31:0] plm_f_data_rsci_q_d_mxwt;
  wire plm_out_data_rsci_bawt;
  wire [31:0] plm_out_data_rsci_q_d_mxwt;
  reg [15:0] dma_read_ctrl_rsci_idat_47_32;
  reg [15:0] dma_read_ctrl_rsci_idat_15_0;
  reg [15:0] dma_write_ctrl_rsci_idat_47_32;
  reg [15:0] dma_write_ctrl_rsci_idat_15_0;
  reg [31:0] dma_write_chnl_rsci_idat_31_0;
  reg CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3;
  reg [29:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4;
  reg CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5;
  wire [3:0] fsm_output;
  wire LOAD_LOOP_LOAD_LOOP_if_and_tmp;
  wire PADDING_LOOP_for_if_equal_tmp;
  wire [8:0] operator_8_false_2_acc_tmp;
  wire [9:0] nl_operator_8_false_2_acc_tmp;
  wire PADDING_LOOP_for_for_if_1_equal_tmp;
  wire [8:0] operator_8_false_1_acc_tmp;
  wire [9:0] nl_operator_8_false_1_acc_tmp;
  wire [5:0] CONVOLUTION_LOOP_acc_tmp;
  wire [6:0] nl_CONVOLUTION_LOOP_acc_tmp;
  wire CONVOLUTION_LOOP_if_equal_tmp;
  wire [8:0] operator_8_false_10_acc_tmp;
  wire [9:0] nl_operator_8_false_10_acc_tmp;
  wire [5:0] CONVOLUTION_LOOP_for_acc_tmp;
  wire [6:0] nl_CONVOLUTION_LOOP_for_acc_tmp;
  wire CONVOLUTION_LOOP_for_for_if_equal_tmp;
  wire [8:0] operator_8_false_8_acc_tmp;
  wire [9:0] nl_operator_8_false_8_acc_tmp;
  wire CONVOLUTION_LOOP_for_for_for_if_2_equal_tmp;
  wire [8:0] operator_8_false_7_acc_tmp;
  wire [9:0] nl_operator_8_false_7_acc_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp;
  wire [8:0] operator_8_false_4_acc_tmp;
  wire [9:0] nl_operator_8_false_4_acc_tmp;
  wire CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_and_1_tmp;
  wire [4:0] BATCH_LOOP_acc_1_tmp;
  wire [5:0] nl_BATCH_LOOP_acc_1_tmp;
  wire BATCH_LOOP_if_2_equal_tmp;
  wire [8:0] operator_8_false_11_acc_tmp;
  wire [9:0] nl_operator_8_false_11_acc_tmp;
  wire STORE_LOOP_if_equal_tmp;
  wire [16:0] operator_16_false_acc_tmp;
  wire [17:0] nl_operator_16_false_acc_tmp;
  wire BATCH_LOOP_and_6_tmp;
  wire STORE_LOOP_STORE_LOOP_or_tmp;
  wire STORE_LOOP_or_2336_tmp;
  wire STORE_LOOP_or_2335_tmp;
  wire BATCH_LOOP_and_4_tmp;
  wire or_tmp_16;
  wire or_tmp_17;
  wire not_tmp_164;
  wire or_tmp_284;
  wire and_dcpl_16;
  wire or_dcpl_28;
  wire and_dcpl_19;
  wire and_dcpl_20;
  wire or_tmp_293;
  wire mux_tmp_319;
  wire and_dcpl_22;
  wire and_dcpl_23;
  wire not_tmp_186;
  wire mux_tmp_321;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_45;
  wire and_dcpl_48;
  wire and_dcpl_55;
  wire and_dcpl_65;
  wire or_tmp_314;
  wire nand_tmp_29;
  wire and_dcpl_69;
  wire and_dcpl_74;
  wire mux_tmp_333;
  wire or_dcpl_48;
  wire or_dcpl_51;
  wire or_tmp_367;
  wire or_tmp_368;
  wire mux_tmp_351;
  wire or_dcpl_56;
  wire or_tmp_369;
  wire mux_tmp_352;
  wire or_tmp_372;
  wire mux_tmp_354;
  wire not_tmp_219;
  wire nand_tmp_39;
  wire mux_tmp_355;
  wire or_dcpl_60;
  wire nor_tmp_142;
  wire mux_tmp_356;
  wire mux_tmp_357;
  wire or_dcpl_65;
  wire and_dcpl_79;
  wire mux_tmp_361;
  wire or_tmp_405;
  wire or_tmp_439;
  wire or_tmp_440;
  wire or_tmp_444;
  wire or_tmp_449;
  wire or_tmp_450;
  wire mux_tmp_372;
  wire or_dcpl_73;
  wire or_tmp_470;
  wire mux_tmp_393;
  wire or_tmp_473;
  wire mux_tmp_395;
  wire or_tmp_492;
  wire or_tmp_496;
  wire mux_tmp_421;
  wire or_tmp_509;
  wire not_tmp_256;
  wire mux_tmp_435;
  wire not_tmp_258;
  wire mux_tmp_446;
  wire mux_tmp_447;
  wire mux_tmp_468;
  wire or_dcpl_85;
  wire or_dcpl_87;
  wire or_dcpl_88;
  wire not_tmp_275;
  wire mux_tmp_472;
  wire not_tmp_291;
  wire and_dcpl_107;
  wire and_dcpl_109;
  wire mux_tmp_510;
  wire or_tmp_625;
  wire mux_tmp_512;
  wire or_tmp_645;
  wire and_dcpl_128;
  wire not_tmp_312;
  wire nand_tmp_57;
  wire and_dcpl_138;
  wire or_dcpl_124;
  wire or_dcpl_127;
  wire and_dcpl_145;
  wire and_dcpl_150;
  wire or_tmp_676;
  wire or_tmp_685;
  wire or_tmp_693;
  wire or_tmp_700;
  wire or_tmp_709;
  wire or_tmp_714;
  wire or_tmp_715;
  wire or_tmp_717;
  wire or_tmp_760;
  wire or_tmp_801;
  wire or_tmp_805;
  wire or_tmp_841;
  wire or_tmp_851;
  wire or_tmp_901;
  wire exit_BATCH_LOOP_sva_2;
  wire exit_STORE_LOOP_lpi_2_dfm_1;
  wire STORE_LOOP_equal_tmp_4;
  wire [15:0] LOAD_LOOP_i_lpi_2_mx1;
  wire [32:0] operator_32_false_acc_psp_sva_1;
  wire [33:0] nl_operator_32_false_acc_psp_sva_1;
  reg [4:0] PADDING_LOOP_chan_5_0_lpi_2_4_0;
  wire exit_PADDING_LOOP_for_for_lpi_2_dfm_1;
  wire exit_PADDING_LOOP_for_sva_5;
  wire exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4;
  wire exit_CONVOLUTION_LOOP_sva_2;
  wire exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4;
  wire exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_sva_5;
  wire CONVOLUTION_LOOP_for_for_for_for_for_if_nor_cse_sva_1;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2;
  reg lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2;
  wire exit_STORE_LOOP_sva_3;
  wire lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0;
  wire lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1;
  wire lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1;
  wire lfst_exit_STORE_LOOP_lpi_2_2_mx1;
  wire lfst_exit_STORE_LOOP_lpi_2_0_mx1;
  wire lfst_exit_STORE_LOOP_lpi_2_1_mx1;
  wire [10:0] buf_acc_data_0_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_0_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_1_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_2_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_3_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_4_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_5_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_6_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_7_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_8_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_9_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_10_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_11_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_12_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_13_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_14_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_15_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_16_17_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_0_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_1_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_2_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_3_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_4_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_5_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_6_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_7_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_8_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_9_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_10_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_11_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_12_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_13_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_14_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_15_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_16_56_46_sva_dfm_1;
  wire [10:0] buf_acc_data_17_17_56_46_sva_dfm_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1;
  reg CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1;
  reg CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0;
  reg [10:0] CONVOLUTION_LOOP_for_for_for_else_mux_itm_1;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1;
  wire CONVOLUTION_LOOP_for_for_for_acc_46_sva_2;
  wire [44:0] CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2;
  wire CONVOLUTION_LOOP_for_for_for_acc_0_sva_2;
  wire [48:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1;
  wire [49:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0;
  reg BATCH_LOOP_stage_v_2;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_2;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_0;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_1;
  reg BATCH_LOOP_stage_v_4;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0;
  reg BATCH_LOOP_stage_v_3;
  wire STORE_LOOP_and_tmp_1;
  wire STORE_LOOP_equal_tmp_6;
  wire STORE_LOOP_equal_tmp_5;
  wire STORE_LOOP_equal_tmp_2_mx0w0;
  wire STORE_LOOP_or_tmp_2;
  reg lfst_exit_PADDING_LOOP_for_lpi_2;
  wire STORE_LOOP_or_tmp_mx0w0;
  reg lfst_exit_CONVOLUTION_LOOP_for_lpi_2;
  wire [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1;
  wire exit_PADDING_LOOP_sva_2;
  wire exit_PADDING_LOOP_for_lpi_2_dfm_4;
  wire [5:0] PADDING_LOOP_chan_5_0_sva_2;
  wire [6:0] nl_PADDING_LOOP_chan_5_0_sva_2;
  reg [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1;
  wire [4:0] CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2;
  reg BATCH_LOOP_asn_itm_1;
  reg exit_BATCH_LOOP_lpi_2_dfm_2_1;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1;
  reg STORE_LOOP_and_35_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1;
  reg BATCH_LOOP_stage_0_4;
  reg BATCH_LOOP_stage_0_2;
  reg BATCH_LOOP_stage_0_3;
  reg lfst_exit_STORE_LOOP_lpi_2_0;
  reg lfst_exit_STORE_LOOP_lpi_2_1;
  reg lfst_exit_STORE_LOOP_lpi_2_2;
  reg exitL_exit_STORE_LOOP_sva;
  reg BATCH_LOOP_stage_0;
  reg STORE_LOOP_equal_tmp_2_1;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_1;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_2;
  reg BATCH_LOOP_asn_itm_2;
  reg STORE_LOOP_equal_tmp_2_2;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2;
  reg BATCH_LOOP_stage_0_1;
  reg lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2;
  reg lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2;
  reg STORE_LOOP_and_15_itm_1;
  reg PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1;
  reg exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1;
  reg [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0;
  reg [4:0] CONVOLUTION_LOOP_for_k_slc_CONVOLUTION_LOOP_for_k_5_0_4_0_3_itm_1;
  reg BATCH_LOOP_stage_v;
  wire exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0;
  reg exit_PADDING_LOOP_for_lpi_2_dfm_1;
  wire exit_CONVOLUTION_LOOP_lpi_2_dfm_mx0w0;
  reg exit_CONVOLUTION_LOOP_lpi_2_dfm;
  wire exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0;
  wire [48:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1;
  wire [49:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1;
  wire exit_LOAD_LOOP_lpi_2_dfm_1;
  wire exit_PADDING_LOOP_lpi_2_dfm_3;
  wire exit_CONVOLUTION_LOOP_lpi_2_dfm_2_mx0w0;
  wire CONVOLUTION_LOOP_for_for_and_psp_mx1w0;
  wire exit_PADDING_LOOP_lpi_2_dfm_mx0w0;
  reg exit_PADDING_LOOP_lpi_2_dfm;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2;
  wire STORE_LOOP_and_11_m1c;
  wire exitL_exit_STORE_LOOP_sva_mx1;
  wire [44:0] CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_45_1_1;
  wire [57:0] CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1;
  wire [58:0] nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1;
  wire [10:0] CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_56_46_1;
  wire STORE_LOOP_and_9_m1c;
  reg reg_CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_ftd_4;
  wire BATCH_LOOP_and_cse;
  wire LOAD_CTRL_LOOP_and_cse;
  reg reg_plm_out_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse;
  reg reg_plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse;
  reg reg_plm_f_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse;
  reg reg_plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse;
  reg reg_plm_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse;
  reg reg_acc_done_rsci_ivld_core_psct_cse;
  reg reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  reg reg_dma_read_chnl_rsci_irdy_core_psct_cse;
  reg reg_dma_write_ctrl_rsci_ivld_core_psct_cse;
  reg reg_dma_read_ctrl_rsci_ivld_core_psct_cse;
  reg reg_conf_info_rsci_irdy_core_psct_cse;
  wire STORE_LOOP_and_703_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_cse;
  wire STORE_LOOP_and_709_cse;
  wire PADDING_LOOP_chan_and_cse;
  wire and_769_cse;
  wire and_770_cse;
  wire nor_240_cse;
  wire and_830_cse;
  wire or_81_cse;
  wire or_214_cse;
  wire BATCH_LOOP_and_10_cse;
  wire PADDING_LOOP_for_for_aelse_2_and_1_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_and_cse;
  wire CONVOLUTION_LOOP_for_for_for_else_and_837_cse;
  wire CONVOLUTION_LOOP_for_for_for_else_and_836_cse;
  wire CONVOLUTION_LOOP_for_for_for_else_and_841_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_and_833_cse;
  wire CONVOLUTION_LOOP_for_for_and_3_cse;
  wire CONVOLUTION_LOOP_for_for_for_acc_and_1_cse;
  wire STORE_LOOP_and_726_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_1_equal_cse;
  wire CONVOLUTION_LOOP_for_if_nor_cse;
  wire or_306_cse;
  wire or_2_cse;
  wire nor_21_cse;
  wire or_1098_cse;
  wire and_831_cse;
  wire nor_229_cse;
  wire nor_93_cse;
  wire nor_90_cse;
  wire nand_109_cse;
  wire or_156_cse;
  wire mux_376_cse;
  wire or_1078_cse;
  wire or_131_cse;
  wire or_1062_cse;
  wire or_141_cse;
  wire or_1096_cse;
  wire or_619_cse;
  wire or_618_cse;
  wire or_617_cse;
  wire or_453_cse;
  wire or_316_cse;
  wire nor_306_cse;
  wire or_668_cse;
  wire nor_303_cse;
  reg STORE_LOOP_or_2332_itm_1;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_2;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_2;
  wire nor_291_cse;
  wire mux_325_cse;
  wire and_765_cse;
  wire or_545_cse;
  wire or_324_cse;
  wire CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_mx0w0;
  wire mux_486_cse;
  wire mux_381_cse_1;
  wire or_548_cse;
  wire mux_490_cse;
  wire mux_484_cse;
  reg [31:0] plm_in_data_rsci_d_d_reg;
  wire [31:0] PADDING_LOOP_for_for_mux_rmff;
  reg [13:0] plm_in_data_rsci_radr_d_reg;
  wire [13:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff;
  reg [13:0] plm_in_data_rsci_wadr_d_reg;
  wire [13:0] PADDING_LOOP_for_for_index_in_mux_rmff;
  wire plm_in_data_rsci_we_d_iff;
  wire and_261_rmff;
  wire plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_253_rmff;
  reg [31:0] plm_f_data_rsci_d_d_reg;
  wire [31:0] LOAD_LOOP_data_ac_mux_rmff;
  reg [15:0] plm_f_data_rsci_radr_d_reg;
  wire [15:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff;
  reg [15:0] plm_f_data_rsci_wadr_d_reg;
  wire [15:0] LOAD_LOOP_i_mux_rmff;
  wire plm_f_data_rsci_we_d_iff;
  wire and_255_rmff;
  wire plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire CONVOLUTION_LOOP_for_for_for_if_1_mux_5_rmff;
  wire [29:0] CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff;
  wire CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff;
  reg [13:0] plm_out_data_rsci_radr_d_reg;
  wire [13:0] CONVOLUTION_LOOP_for_for_for_index_out_mux_1_rmff;
  reg [13:0] plm_out_data_rsci_wadr_d_reg;
  wire [13:0] CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff;
  wire plm_out_data_rsci_we_d_iff;
  wire and_247_rmff;
  wire plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_245_rmff;
  wire and_257_rmff;
  wire or_dcpl_135;
  wire or_dcpl_162;
  wire or_dcpl_163;
  wire or_dcpl_168;
  wire or_dcpl_169;
  wire STORE_LOOP_and_32_cse;
  wire STORE_LOOP_and_4_cse;
  wire STORE_LOOP_and_30_cse;
  wire STORE_LOOP_and_10_cse;
  wire STORE_LOOP_and_12_cse;
  wire [54:0] CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0;
  wire PADDING_LOOP_for_and_tmp_1;
  wire CONVOLUTION_LOOP_for_and_tmp_1;
  reg STORE_LOOP_or_tmp_1;
  reg STORE_LOOP_or_2_itm_1;
  wire PADDING_LOOP_for_for_and_psp_mx1w0;
  wire STORE_LOOP_asn_3330;
  wire STORE_LOOP_and_1_m1c_1;
  wire nor_385_m1c;
  wire nor_384_m1c;
  wire or_1160_tmp;
  wire STORE_LOOP_and_27_tmp;
  wire or_1156_tmp;
  wire and_876_tmp;
  wire STORE_LOOP_and_6_tmp;
  wire or_1135_tmp;
  wire or_1127_tmp;
  wire STORE_LOOP_and_24_tmp;
  wire or_1123_tmp;
  wire STORE_LOOP_and_22_tmp;
  wire STORE_LOOP_and_33_cse;
  wire STORE_LOOP_and_29_cse;
  wire STORE_LOOP_and_31_cse;
  wire or_1066_cse;
  wire or_1067_cse;
  reg CONVOLUTION_LOOP_for_for_and_psp;
  reg PADDING_LOOP_for_for_and_psp;
  wire dma_read_info_index_and_itm;
  wire [15:0] z_out;
  wire [16:0] nl_z_out;
  wire [9:0] z_out_2;
  wire [8:0] z_out_3;
  wire [8:0] z_out_4;
  wire [9:0] nl_z_out_4;
  wire [15:0] z_out_6;
  wire [23:0] nl_z_out_6;
  wire [63:0] z_out_7;
  wire [31:0] z_out_10;
  wire [16:0] z_out_12;
  wire [17:0] nl_z_out_12;
  wire [7:0] z_out_13;
  wire [8:0] nl_z_out_13;
  reg [15:0] dma_read_info_index_15_0_lpi_2;
  reg [15:0] LOAD_LOOP_i_lpi_2;
  reg [4:0] PADDING_LOOP_for_row_4_0_lpi_2;
  reg [4:0] PADDING_LOOP_for_for_col_4_0_lpi_2;
  reg [4:0] CONVOLUTION_LOOP_for_for_i_4_0_lpi_2;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2;
  reg CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2;
  reg CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_2;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_y_lpi_2;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2;
  reg [13:0] STORE_LOOP_i_13_0_lpi_2;
  reg [44:0] buf_acc_data_8_17_45_1_sva;
  reg buf_acc_data_8_17_0_sva;
  reg [10:0] buf_acc_data_8_17_56_46_sva;
  reg [44:0] buf_acc_data_9_0_45_1_sva;
  reg buf_acc_data_9_0_0_sva;
  reg [10:0] buf_acc_data_9_0_56_46_sva;
  reg [44:0] buf_acc_data_8_16_45_1_sva;
  reg buf_acc_data_8_16_0_sva;
  reg [10:0] buf_acc_data_8_16_56_46_sva;
  reg [44:0] buf_acc_data_9_1_45_1_sva;
  reg buf_acc_data_9_1_0_sva;
  reg [10:0] buf_acc_data_9_1_56_46_sva;
  reg [44:0] buf_acc_data_8_15_45_1_sva;
  reg buf_acc_data_8_15_0_sva;
  reg [10:0] buf_acc_data_8_15_56_46_sva;
  reg [44:0] buf_acc_data_9_2_45_1_sva;
  reg buf_acc_data_9_2_0_sva;
  reg [10:0] buf_acc_data_9_2_56_46_sva;
  reg [44:0] buf_acc_data_8_14_45_1_sva;
  reg buf_acc_data_8_14_0_sva;
  reg [10:0] buf_acc_data_8_14_56_46_sva;
  reg [44:0] buf_acc_data_9_3_45_1_sva;
  reg buf_acc_data_9_3_0_sva;
  reg [10:0] buf_acc_data_9_3_56_46_sva;
  reg [44:0] buf_acc_data_8_13_45_1_sva;
  reg buf_acc_data_8_13_0_sva;
  reg [10:0] buf_acc_data_8_13_56_46_sva;
  reg [44:0] buf_acc_data_9_4_45_1_sva;
  reg buf_acc_data_9_4_0_sva;
  reg [10:0] buf_acc_data_9_4_56_46_sva;
  reg [44:0] buf_acc_data_8_12_45_1_sva;
  reg buf_acc_data_8_12_0_sva;
  reg [10:0] buf_acc_data_8_12_56_46_sva;
  reg [44:0] buf_acc_data_9_5_45_1_sva;
  reg buf_acc_data_9_5_0_sva;
  reg [10:0] buf_acc_data_9_5_56_46_sva;
  reg [44:0] buf_acc_data_8_11_45_1_sva;
  reg buf_acc_data_8_11_0_sva;
  reg [10:0] buf_acc_data_8_11_56_46_sva;
  reg [44:0] buf_acc_data_9_6_45_1_sva;
  reg buf_acc_data_9_6_0_sva;
  reg [10:0] buf_acc_data_9_6_56_46_sva;
  reg [44:0] buf_acc_data_8_10_45_1_sva;
  reg buf_acc_data_8_10_0_sva;
  reg [10:0] buf_acc_data_8_10_56_46_sva;
  reg [44:0] buf_acc_data_9_7_45_1_sva;
  reg buf_acc_data_9_7_0_sva;
  reg [10:0] buf_acc_data_9_7_56_46_sva;
  reg [44:0] buf_acc_data_8_9_45_1_sva;
  reg buf_acc_data_8_9_0_sva;
  reg [10:0] buf_acc_data_8_9_56_46_sva;
  reg [44:0] buf_acc_data_9_8_45_1_sva;
  reg buf_acc_data_9_8_0_sva;
  reg [10:0] buf_acc_data_9_8_56_46_sva;
  reg [44:0] buf_acc_data_8_8_45_1_sva;
  reg buf_acc_data_8_8_0_sva;
  reg [10:0] buf_acc_data_8_8_56_46_sva;
  reg [44:0] buf_acc_data_9_9_45_1_sva;
  reg buf_acc_data_9_9_0_sva;
  reg [10:0] buf_acc_data_9_9_56_46_sva;
  reg [44:0] buf_acc_data_8_7_45_1_sva;
  reg buf_acc_data_8_7_0_sva;
  reg [10:0] buf_acc_data_8_7_56_46_sva;
  reg [44:0] buf_acc_data_9_10_45_1_sva;
  reg buf_acc_data_9_10_0_sva;
  reg [10:0] buf_acc_data_9_10_56_46_sva;
  reg [44:0] buf_acc_data_8_6_45_1_sva;
  reg buf_acc_data_8_6_0_sva;
  reg [10:0] buf_acc_data_8_6_56_46_sva;
  reg [44:0] buf_acc_data_9_11_45_1_sva;
  reg buf_acc_data_9_11_0_sva;
  reg [10:0] buf_acc_data_9_11_56_46_sva;
  reg [44:0] buf_acc_data_8_5_45_1_sva;
  reg buf_acc_data_8_5_0_sva;
  reg [10:0] buf_acc_data_8_5_56_46_sva;
  reg [44:0] buf_acc_data_9_12_45_1_sva;
  reg buf_acc_data_9_12_0_sva;
  reg [10:0] buf_acc_data_9_12_56_46_sva;
  reg [44:0] buf_acc_data_8_4_45_1_sva;
  reg buf_acc_data_8_4_0_sva;
  reg [10:0] buf_acc_data_8_4_56_46_sva;
  reg [44:0] buf_acc_data_9_13_45_1_sva;
  reg buf_acc_data_9_13_0_sva;
  reg [10:0] buf_acc_data_9_13_56_46_sva;
  reg [44:0] buf_acc_data_8_3_45_1_sva;
  reg buf_acc_data_8_3_0_sva;
  reg [10:0] buf_acc_data_8_3_56_46_sva;
  reg [44:0] buf_acc_data_9_14_45_1_sva;
  reg buf_acc_data_9_14_0_sva;
  reg [10:0] buf_acc_data_9_14_56_46_sva;
  reg [44:0] buf_acc_data_8_2_45_1_sva;
  reg buf_acc_data_8_2_0_sva;
  reg [10:0] buf_acc_data_8_2_56_46_sva;
  reg [44:0] buf_acc_data_9_15_45_1_sva;
  reg buf_acc_data_9_15_0_sva;
  reg [10:0] buf_acc_data_9_15_56_46_sva;
  reg [44:0] buf_acc_data_8_1_45_1_sva;
  reg buf_acc_data_8_1_0_sva;
  reg [10:0] buf_acc_data_8_1_56_46_sva;
  reg [44:0] buf_acc_data_9_16_45_1_sva;
  reg buf_acc_data_9_16_0_sva;
  reg [10:0] buf_acc_data_9_16_56_46_sva;
  reg [44:0] buf_acc_data_8_0_45_1_sva;
  reg buf_acc_data_8_0_0_sva;
  reg [10:0] buf_acc_data_8_0_56_46_sva;
  reg [44:0] buf_acc_data_9_17_45_1_sva;
  reg buf_acc_data_9_17_0_sva;
  reg [10:0] buf_acc_data_9_17_56_46_sva;
  reg [44:0] buf_acc_data_7_17_45_1_sva;
  reg buf_acc_data_7_17_0_sva;
  reg [10:0] buf_acc_data_7_17_56_46_sva;
  reg [44:0] buf_acc_data_10_0_45_1_sva;
  reg buf_acc_data_10_0_0_sva;
  reg [10:0] buf_acc_data_10_0_56_46_sva;
  reg [44:0] buf_acc_data_7_16_45_1_sva;
  reg buf_acc_data_7_16_0_sva;
  reg [10:0] buf_acc_data_7_16_56_46_sva;
  reg [44:0] buf_acc_data_10_1_45_1_sva;
  reg buf_acc_data_10_1_0_sva;
  reg [10:0] buf_acc_data_10_1_56_46_sva;
  reg [44:0] buf_acc_data_7_15_45_1_sva;
  reg buf_acc_data_7_15_0_sva;
  reg [10:0] buf_acc_data_7_15_56_46_sva;
  reg [44:0] buf_acc_data_10_2_45_1_sva;
  reg buf_acc_data_10_2_0_sva;
  reg [10:0] buf_acc_data_10_2_56_46_sva;
  reg [44:0] buf_acc_data_7_14_45_1_sva;
  reg buf_acc_data_7_14_0_sva;
  reg [10:0] buf_acc_data_7_14_56_46_sva;
  reg [44:0] buf_acc_data_10_3_45_1_sva;
  reg buf_acc_data_10_3_0_sva;
  reg [10:0] buf_acc_data_10_3_56_46_sva;
  reg [44:0] buf_acc_data_7_13_45_1_sva;
  reg buf_acc_data_7_13_0_sva;
  reg [10:0] buf_acc_data_7_13_56_46_sva;
  reg [44:0] buf_acc_data_10_4_45_1_sva;
  reg buf_acc_data_10_4_0_sva;
  reg [10:0] buf_acc_data_10_4_56_46_sva;
  reg [44:0] buf_acc_data_7_12_45_1_sva;
  reg buf_acc_data_7_12_0_sva;
  reg [10:0] buf_acc_data_7_12_56_46_sva;
  reg [44:0] buf_acc_data_10_5_45_1_sva;
  reg buf_acc_data_10_5_0_sva;
  reg [10:0] buf_acc_data_10_5_56_46_sva;
  reg [44:0] buf_acc_data_7_11_45_1_sva;
  reg buf_acc_data_7_11_0_sva;
  reg [10:0] buf_acc_data_7_11_56_46_sva;
  reg [44:0] buf_acc_data_10_6_45_1_sva;
  reg buf_acc_data_10_6_0_sva;
  reg [10:0] buf_acc_data_10_6_56_46_sva;
  reg [44:0] buf_acc_data_7_10_45_1_sva;
  reg buf_acc_data_7_10_0_sva;
  reg [10:0] buf_acc_data_7_10_56_46_sva;
  reg [44:0] buf_acc_data_10_7_45_1_sva;
  reg buf_acc_data_10_7_0_sva;
  reg [10:0] buf_acc_data_10_7_56_46_sva;
  reg [44:0] buf_acc_data_7_9_45_1_sva;
  reg buf_acc_data_7_9_0_sva;
  reg [10:0] buf_acc_data_7_9_56_46_sva;
  reg [44:0] buf_acc_data_10_8_45_1_sva;
  reg buf_acc_data_10_8_0_sva;
  reg [10:0] buf_acc_data_10_8_56_46_sva;
  reg [44:0] buf_acc_data_7_8_45_1_sva;
  reg buf_acc_data_7_8_0_sva;
  reg [10:0] buf_acc_data_7_8_56_46_sva;
  reg [44:0] buf_acc_data_10_9_45_1_sva;
  reg buf_acc_data_10_9_0_sva;
  reg [10:0] buf_acc_data_10_9_56_46_sva;
  reg [44:0] buf_acc_data_7_7_45_1_sva;
  reg buf_acc_data_7_7_0_sva;
  reg [10:0] buf_acc_data_7_7_56_46_sva;
  reg [44:0] buf_acc_data_10_10_45_1_sva;
  reg buf_acc_data_10_10_0_sva;
  reg [10:0] buf_acc_data_10_10_56_46_sva;
  reg [44:0] buf_acc_data_7_6_45_1_sva;
  reg buf_acc_data_7_6_0_sva;
  reg [10:0] buf_acc_data_7_6_56_46_sva;
  reg [44:0] buf_acc_data_10_11_45_1_sva;
  reg buf_acc_data_10_11_0_sva;
  reg [10:0] buf_acc_data_10_11_56_46_sva;
  reg [44:0] buf_acc_data_7_5_45_1_sva;
  reg buf_acc_data_7_5_0_sva;
  reg [10:0] buf_acc_data_7_5_56_46_sva;
  reg [44:0] buf_acc_data_10_12_45_1_sva;
  reg buf_acc_data_10_12_0_sva;
  reg [10:0] buf_acc_data_10_12_56_46_sva;
  reg [44:0] buf_acc_data_7_4_45_1_sva;
  reg buf_acc_data_7_4_0_sva;
  reg [10:0] buf_acc_data_7_4_56_46_sva;
  reg [44:0] buf_acc_data_10_13_45_1_sva;
  reg buf_acc_data_10_13_0_sva;
  reg [10:0] buf_acc_data_10_13_56_46_sva;
  reg [44:0] buf_acc_data_7_3_45_1_sva;
  reg buf_acc_data_7_3_0_sva;
  reg [10:0] buf_acc_data_7_3_56_46_sva;
  reg [44:0] buf_acc_data_10_14_45_1_sva;
  reg buf_acc_data_10_14_0_sva;
  reg [10:0] buf_acc_data_10_14_56_46_sva;
  reg [44:0] buf_acc_data_7_2_45_1_sva;
  reg buf_acc_data_7_2_0_sva;
  reg [10:0] buf_acc_data_7_2_56_46_sva;
  reg [44:0] buf_acc_data_10_15_45_1_sva;
  reg buf_acc_data_10_15_0_sva;
  reg [10:0] buf_acc_data_10_15_56_46_sva;
  reg [44:0] buf_acc_data_7_1_45_1_sva;
  reg buf_acc_data_7_1_0_sva;
  reg [10:0] buf_acc_data_7_1_56_46_sva;
  reg [44:0] buf_acc_data_10_16_45_1_sva;
  reg buf_acc_data_10_16_0_sva;
  reg [10:0] buf_acc_data_10_16_56_46_sva;
  reg [44:0] buf_acc_data_7_0_45_1_sva;
  reg buf_acc_data_7_0_0_sva;
  reg [10:0] buf_acc_data_7_0_56_46_sva;
  reg [44:0] buf_acc_data_10_17_45_1_sva;
  reg buf_acc_data_10_17_0_sva;
  reg [10:0] buf_acc_data_10_17_56_46_sva;
  reg [44:0] buf_acc_data_6_17_45_1_sva;
  reg buf_acc_data_6_17_0_sva;
  reg [10:0] buf_acc_data_6_17_56_46_sva;
  reg [44:0] buf_acc_data_11_0_45_1_sva;
  reg buf_acc_data_11_0_0_sva;
  reg [10:0] buf_acc_data_11_0_56_46_sva;
  reg [44:0] buf_acc_data_6_16_45_1_sva;
  reg buf_acc_data_6_16_0_sva;
  reg [10:0] buf_acc_data_6_16_56_46_sva;
  reg [44:0] buf_acc_data_11_1_45_1_sva;
  reg buf_acc_data_11_1_0_sva;
  reg [10:0] buf_acc_data_11_1_56_46_sva;
  reg [44:0] buf_acc_data_6_15_45_1_sva;
  reg buf_acc_data_6_15_0_sva;
  reg [10:0] buf_acc_data_6_15_56_46_sva;
  reg [44:0] buf_acc_data_11_2_45_1_sva;
  reg buf_acc_data_11_2_0_sva;
  reg [10:0] buf_acc_data_11_2_56_46_sva;
  reg [44:0] buf_acc_data_6_14_45_1_sva;
  reg buf_acc_data_6_14_0_sva;
  reg [10:0] buf_acc_data_6_14_56_46_sva;
  reg [44:0] buf_acc_data_11_3_45_1_sva;
  reg buf_acc_data_11_3_0_sva;
  reg [10:0] buf_acc_data_11_3_56_46_sva;
  reg [44:0] buf_acc_data_6_13_45_1_sva;
  reg buf_acc_data_6_13_0_sva;
  reg [10:0] buf_acc_data_6_13_56_46_sva;
  reg [44:0] buf_acc_data_11_4_45_1_sva;
  reg buf_acc_data_11_4_0_sva;
  reg [10:0] buf_acc_data_11_4_56_46_sva;
  reg [44:0] buf_acc_data_6_12_45_1_sva;
  reg buf_acc_data_6_12_0_sva;
  reg [10:0] buf_acc_data_6_12_56_46_sva;
  reg [44:0] buf_acc_data_11_5_45_1_sva;
  reg buf_acc_data_11_5_0_sva;
  reg [10:0] buf_acc_data_11_5_56_46_sva;
  reg [44:0] buf_acc_data_6_11_45_1_sva;
  reg buf_acc_data_6_11_0_sva;
  reg [10:0] buf_acc_data_6_11_56_46_sva;
  reg [44:0] buf_acc_data_11_6_45_1_sva;
  reg buf_acc_data_11_6_0_sva;
  reg [10:0] buf_acc_data_11_6_56_46_sva;
  reg [44:0] buf_acc_data_6_10_45_1_sva;
  reg buf_acc_data_6_10_0_sva;
  reg [10:0] buf_acc_data_6_10_56_46_sva;
  reg [44:0] buf_acc_data_11_7_45_1_sva;
  reg buf_acc_data_11_7_0_sva;
  reg [10:0] buf_acc_data_11_7_56_46_sva;
  reg [44:0] buf_acc_data_6_9_45_1_sva;
  reg buf_acc_data_6_9_0_sva;
  reg [10:0] buf_acc_data_6_9_56_46_sva;
  reg [44:0] buf_acc_data_11_8_45_1_sva;
  reg buf_acc_data_11_8_0_sva;
  reg [10:0] buf_acc_data_11_8_56_46_sva;
  reg [44:0] buf_acc_data_6_8_45_1_sva;
  reg buf_acc_data_6_8_0_sva;
  reg [10:0] buf_acc_data_6_8_56_46_sva;
  reg [44:0] buf_acc_data_11_9_45_1_sva;
  reg buf_acc_data_11_9_0_sva;
  reg [10:0] buf_acc_data_11_9_56_46_sva;
  reg [44:0] buf_acc_data_6_7_45_1_sva;
  reg buf_acc_data_6_7_0_sva;
  reg [10:0] buf_acc_data_6_7_56_46_sva;
  reg [44:0] buf_acc_data_11_10_45_1_sva;
  reg buf_acc_data_11_10_0_sva;
  reg [10:0] buf_acc_data_11_10_56_46_sva;
  reg [44:0] buf_acc_data_6_6_45_1_sva;
  reg buf_acc_data_6_6_0_sva;
  reg [10:0] buf_acc_data_6_6_56_46_sva;
  reg [44:0] buf_acc_data_11_11_45_1_sva;
  reg buf_acc_data_11_11_0_sva;
  reg [10:0] buf_acc_data_11_11_56_46_sva;
  reg [44:0] buf_acc_data_6_5_45_1_sva;
  reg buf_acc_data_6_5_0_sva;
  reg [10:0] buf_acc_data_6_5_56_46_sva;
  reg [44:0] buf_acc_data_11_12_45_1_sva;
  reg buf_acc_data_11_12_0_sva;
  reg [10:0] buf_acc_data_11_12_56_46_sva;
  reg [44:0] buf_acc_data_6_4_45_1_sva;
  reg buf_acc_data_6_4_0_sva;
  reg [10:0] buf_acc_data_6_4_56_46_sva;
  reg [44:0] buf_acc_data_11_13_45_1_sva;
  reg buf_acc_data_11_13_0_sva;
  reg [10:0] buf_acc_data_11_13_56_46_sva;
  reg [44:0] buf_acc_data_6_3_45_1_sva;
  reg buf_acc_data_6_3_0_sva;
  reg [10:0] buf_acc_data_6_3_56_46_sva;
  reg [44:0] buf_acc_data_11_14_45_1_sva;
  reg buf_acc_data_11_14_0_sva;
  reg [10:0] buf_acc_data_11_14_56_46_sva;
  reg [44:0] buf_acc_data_6_2_45_1_sva;
  reg buf_acc_data_6_2_0_sva;
  reg [10:0] buf_acc_data_6_2_56_46_sva;
  reg [44:0] buf_acc_data_11_15_45_1_sva;
  reg buf_acc_data_11_15_0_sva;
  reg [10:0] buf_acc_data_11_15_56_46_sva;
  reg [44:0] buf_acc_data_6_1_45_1_sva;
  reg buf_acc_data_6_1_0_sva;
  reg [10:0] buf_acc_data_6_1_56_46_sva;
  reg [44:0] buf_acc_data_11_16_45_1_sva;
  reg buf_acc_data_11_16_0_sva;
  reg [10:0] buf_acc_data_11_16_56_46_sva;
  reg [44:0] buf_acc_data_6_0_45_1_sva;
  reg buf_acc_data_6_0_0_sva;
  reg [10:0] buf_acc_data_6_0_56_46_sva;
  reg [44:0] buf_acc_data_11_17_45_1_sva;
  reg buf_acc_data_11_17_0_sva;
  reg [10:0] buf_acc_data_11_17_56_46_sva;
  reg [44:0] buf_acc_data_5_17_45_1_sva;
  reg buf_acc_data_5_17_0_sva;
  reg [10:0] buf_acc_data_5_17_56_46_sva;
  reg [44:0] buf_acc_data_12_0_45_1_sva;
  reg buf_acc_data_12_0_0_sva;
  reg [10:0] buf_acc_data_12_0_56_46_sva;
  reg [44:0] buf_acc_data_5_16_45_1_sva;
  reg buf_acc_data_5_16_0_sva;
  reg [10:0] buf_acc_data_5_16_56_46_sva;
  reg [44:0] buf_acc_data_12_1_45_1_sva;
  reg buf_acc_data_12_1_0_sva;
  reg [10:0] buf_acc_data_12_1_56_46_sva;
  reg [44:0] buf_acc_data_5_15_45_1_sva;
  reg buf_acc_data_5_15_0_sva;
  reg [10:0] buf_acc_data_5_15_56_46_sva;
  reg [44:0] buf_acc_data_12_2_45_1_sva;
  reg buf_acc_data_12_2_0_sva;
  reg [10:0] buf_acc_data_12_2_56_46_sva;
  reg [44:0] buf_acc_data_5_14_45_1_sva;
  reg buf_acc_data_5_14_0_sva;
  reg [10:0] buf_acc_data_5_14_56_46_sva;
  reg [44:0] buf_acc_data_12_3_45_1_sva;
  reg buf_acc_data_12_3_0_sva;
  reg [10:0] buf_acc_data_12_3_56_46_sva;
  reg [44:0] buf_acc_data_5_13_45_1_sva;
  reg buf_acc_data_5_13_0_sva;
  reg [10:0] buf_acc_data_5_13_56_46_sva;
  reg [44:0] buf_acc_data_12_4_45_1_sva;
  reg buf_acc_data_12_4_0_sva;
  reg [10:0] buf_acc_data_12_4_56_46_sva;
  reg [44:0] buf_acc_data_5_12_45_1_sva;
  reg buf_acc_data_5_12_0_sva;
  reg [10:0] buf_acc_data_5_12_56_46_sva;
  reg [44:0] buf_acc_data_12_5_45_1_sva;
  reg buf_acc_data_12_5_0_sva;
  reg [10:0] buf_acc_data_12_5_56_46_sva;
  reg [44:0] buf_acc_data_5_11_45_1_sva;
  reg buf_acc_data_5_11_0_sva;
  reg [10:0] buf_acc_data_5_11_56_46_sva;
  reg [44:0] buf_acc_data_12_6_45_1_sva;
  reg buf_acc_data_12_6_0_sva;
  reg [10:0] buf_acc_data_12_6_56_46_sva;
  reg [44:0] buf_acc_data_5_10_45_1_sva;
  reg buf_acc_data_5_10_0_sva;
  reg [10:0] buf_acc_data_5_10_56_46_sva;
  reg [44:0] buf_acc_data_12_7_45_1_sva;
  reg buf_acc_data_12_7_0_sva;
  reg [10:0] buf_acc_data_12_7_56_46_sva;
  reg [44:0] buf_acc_data_5_9_45_1_sva;
  reg buf_acc_data_5_9_0_sva;
  reg [10:0] buf_acc_data_5_9_56_46_sva;
  reg [44:0] buf_acc_data_12_8_45_1_sva;
  reg buf_acc_data_12_8_0_sva;
  reg [10:0] buf_acc_data_12_8_56_46_sva;
  reg [44:0] buf_acc_data_5_8_45_1_sva;
  reg buf_acc_data_5_8_0_sva;
  reg [10:0] buf_acc_data_5_8_56_46_sva;
  reg [44:0] buf_acc_data_12_9_45_1_sva;
  reg buf_acc_data_12_9_0_sva;
  reg [10:0] buf_acc_data_12_9_56_46_sva;
  reg [44:0] buf_acc_data_5_7_45_1_sva;
  reg buf_acc_data_5_7_0_sva;
  reg [10:0] buf_acc_data_5_7_56_46_sva;
  reg [44:0] buf_acc_data_12_10_45_1_sva;
  reg buf_acc_data_12_10_0_sva;
  reg [10:0] buf_acc_data_12_10_56_46_sva;
  reg [44:0] buf_acc_data_5_6_45_1_sva;
  reg buf_acc_data_5_6_0_sva;
  reg [10:0] buf_acc_data_5_6_56_46_sva;
  reg [44:0] buf_acc_data_12_11_45_1_sva;
  reg buf_acc_data_12_11_0_sva;
  reg [10:0] buf_acc_data_12_11_56_46_sva;
  reg [44:0] buf_acc_data_5_5_45_1_sva;
  reg buf_acc_data_5_5_0_sva;
  reg [10:0] buf_acc_data_5_5_56_46_sva;
  reg [44:0] buf_acc_data_12_12_45_1_sva;
  reg buf_acc_data_12_12_0_sva;
  reg [10:0] buf_acc_data_12_12_56_46_sva;
  reg [44:0] buf_acc_data_5_4_45_1_sva;
  reg buf_acc_data_5_4_0_sva;
  reg [10:0] buf_acc_data_5_4_56_46_sva;
  reg [44:0] buf_acc_data_12_13_45_1_sva;
  reg buf_acc_data_12_13_0_sva;
  reg [10:0] buf_acc_data_12_13_56_46_sva;
  reg [44:0] buf_acc_data_5_3_45_1_sva;
  reg buf_acc_data_5_3_0_sva;
  reg [10:0] buf_acc_data_5_3_56_46_sva;
  reg [44:0] buf_acc_data_12_14_45_1_sva;
  reg buf_acc_data_12_14_0_sva;
  reg [10:0] buf_acc_data_12_14_56_46_sva;
  reg [44:0] buf_acc_data_5_2_45_1_sva;
  reg buf_acc_data_5_2_0_sva;
  reg [10:0] buf_acc_data_5_2_56_46_sva;
  reg [44:0] buf_acc_data_12_15_45_1_sva;
  reg buf_acc_data_12_15_0_sva;
  reg [10:0] buf_acc_data_12_15_56_46_sva;
  reg [44:0] buf_acc_data_5_1_45_1_sva;
  reg buf_acc_data_5_1_0_sva;
  reg [10:0] buf_acc_data_5_1_56_46_sva;
  reg [44:0] buf_acc_data_12_16_45_1_sva;
  reg buf_acc_data_12_16_0_sva;
  reg [10:0] buf_acc_data_12_16_56_46_sva;
  reg [44:0] buf_acc_data_5_0_45_1_sva;
  reg buf_acc_data_5_0_0_sva;
  reg [10:0] buf_acc_data_5_0_56_46_sva;
  reg [44:0] buf_acc_data_12_17_45_1_sva;
  reg buf_acc_data_12_17_0_sva;
  reg [10:0] buf_acc_data_12_17_56_46_sva;
  reg [44:0] buf_acc_data_4_17_45_1_sva;
  reg buf_acc_data_4_17_0_sva;
  reg [10:0] buf_acc_data_4_17_56_46_sva;
  reg [44:0] buf_acc_data_13_0_45_1_sva;
  reg buf_acc_data_13_0_0_sva;
  reg [10:0] buf_acc_data_13_0_56_46_sva;
  reg [44:0] buf_acc_data_4_16_45_1_sva;
  reg buf_acc_data_4_16_0_sva;
  reg [10:0] buf_acc_data_4_16_56_46_sva;
  reg [44:0] buf_acc_data_13_1_45_1_sva;
  reg buf_acc_data_13_1_0_sva;
  reg [10:0] buf_acc_data_13_1_56_46_sva;
  reg [44:0] buf_acc_data_4_15_45_1_sva;
  reg buf_acc_data_4_15_0_sva;
  reg [10:0] buf_acc_data_4_15_56_46_sva;
  reg [44:0] buf_acc_data_13_2_45_1_sva;
  reg buf_acc_data_13_2_0_sva;
  reg [10:0] buf_acc_data_13_2_56_46_sva;
  reg [44:0] buf_acc_data_4_14_45_1_sva;
  reg buf_acc_data_4_14_0_sva;
  reg [10:0] buf_acc_data_4_14_56_46_sva;
  reg [44:0] buf_acc_data_13_3_45_1_sva;
  reg buf_acc_data_13_3_0_sva;
  reg [10:0] buf_acc_data_13_3_56_46_sva;
  reg [44:0] buf_acc_data_4_13_45_1_sva;
  reg buf_acc_data_4_13_0_sva;
  reg [10:0] buf_acc_data_4_13_56_46_sva;
  reg [44:0] buf_acc_data_13_4_45_1_sva;
  reg buf_acc_data_13_4_0_sva;
  reg [10:0] buf_acc_data_13_4_56_46_sva;
  reg [44:0] buf_acc_data_4_12_45_1_sva;
  reg buf_acc_data_4_12_0_sva;
  reg [10:0] buf_acc_data_4_12_56_46_sva;
  reg [44:0] buf_acc_data_13_5_45_1_sva;
  reg buf_acc_data_13_5_0_sva;
  reg [10:0] buf_acc_data_13_5_56_46_sva;
  reg [44:0] buf_acc_data_4_11_45_1_sva;
  reg buf_acc_data_4_11_0_sva;
  reg [10:0] buf_acc_data_4_11_56_46_sva;
  reg [44:0] buf_acc_data_13_6_45_1_sva;
  reg buf_acc_data_13_6_0_sva;
  reg [10:0] buf_acc_data_13_6_56_46_sva;
  reg [44:0] buf_acc_data_4_10_45_1_sva;
  reg buf_acc_data_4_10_0_sva;
  reg [10:0] buf_acc_data_4_10_56_46_sva;
  reg [44:0] buf_acc_data_13_7_45_1_sva;
  reg buf_acc_data_13_7_0_sva;
  reg [10:0] buf_acc_data_13_7_56_46_sva;
  reg [44:0] buf_acc_data_4_9_45_1_sva;
  reg buf_acc_data_4_9_0_sva;
  reg [10:0] buf_acc_data_4_9_56_46_sva;
  reg [44:0] buf_acc_data_13_8_45_1_sva;
  reg buf_acc_data_13_8_0_sva;
  reg [10:0] buf_acc_data_13_8_56_46_sva;
  reg [44:0] buf_acc_data_4_8_45_1_sva;
  reg buf_acc_data_4_8_0_sva;
  reg [10:0] buf_acc_data_4_8_56_46_sva;
  reg [44:0] buf_acc_data_13_9_45_1_sva;
  reg buf_acc_data_13_9_0_sva;
  reg [10:0] buf_acc_data_13_9_56_46_sva;
  reg [44:0] buf_acc_data_4_7_45_1_sva;
  reg buf_acc_data_4_7_0_sva;
  reg [10:0] buf_acc_data_4_7_56_46_sva;
  reg [44:0] buf_acc_data_13_10_45_1_sva;
  reg buf_acc_data_13_10_0_sva;
  reg [10:0] buf_acc_data_13_10_56_46_sva;
  reg [44:0] buf_acc_data_4_6_45_1_sva;
  reg buf_acc_data_4_6_0_sva;
  reg [10:0] buf_acc_data_4_6_56_46_sva;
  reg [44:0] buf_acc_data_13_11_45_1_sva;
  reg buf_acc_data_13_11_0_sva;
  reg [10:0] buf_acc_data_13_11_56_46_sva;
  reg [44:0] buf_acc_data_4_5_45_1_sva;
  reg buf_acc_data_4_5_0_sva;
  reg [10:0] buf_acc_data_4_5_56_46_sva;
  reg [44:0] buf_acc_data_13_12_45_1_sva;
  reg buf_acc_data_13_12_0_sva;
  reg [10:0] buf_acc_data_13_12_56_46_sva;
  reg [44:0] buf_acc_data_4_4_45_1_sva;
  reg buf_acc_data_4_4_0_sva;
  reg [10:0] buf_acc_data_4_4_56_46_sva;
  reg [44:0] buf_acc_data_13_13_45_1_sva;
  reg buf_acc_data_13_13_0_sva;
  reg [10:0] buf_acc_data_13_13_56_46_sva;
  reg [44:0] buf_acc_data_4_3_45_1_sva;
  reg buf_acc_data_4_3_0_sva;
  reg [10:0] buf_acc_data_4_3_56_46_sva;
  reg [44:0] buf_acc_data_13_14_45_1_sva;
  reg buf_acc_data_13_14_0_sva;
  reg [10:0] buf_acc_data_13_14_56_46_sva;
  reg [44:0] buf_acc_data_4_2_45_1_sva;
  reg buf_acc_data_4_2_0_sva;
  reg [10:0] buf_acc_data_4_2_56_46_sva;
  reg [44:0] buf_acc_data_13_15_45_1_sva;
  reg buf_acc_data_13_15_0_sva;
  reg [10:0] buf_acc_data_13_15_56_46_sva;
  reg [44:0] buf_acc_data_4_1_45_1_sva;
  reg buf_acc_data_4_1_0_sva;
  reg [10:0] buf_acc_data_4_1_56_46_sva;
  reg [44:0] buf_acc_data_13_16_45_1_sva;
  reg buf_acc_data_13_16_0_sva;
  reg [10:0] buf_acc_data_13_16_56_46_sva;
  reg [44:0] buf_acc_data_4_0_45_1_sva;
  reg buf_acc_data_4_0_0_sva;
  reg [10:0] buf_acc_data_4_0_56_46_sva;
  reg [44:0] buf_acc_data_13_17_45_1_sva;
  reg buf_acc_data_13_17_0_sva;
  reg [10:0] buf_acc_data_13_17_56_46_sva;
  reg [44:0] buf_acc_data_3_17_45_1_sva;
  reg buf_acc_data_3_17_0_sva;
  reg [10:0] buf_acc_data_3_17_56_46_sva;
  reg [44:0] buf_acc_data_14_0_45_1_sva;
  reg buf_acc_data_14_0_0_sva;
  reg [10:0] buf_acc_data_14_0_56_46_sva;
  reg [44:0] buf_acc_data_3_16_45_1_sva;
  reg buf_acc_data_3_16_0_sva;
  reg [10:0] buf_acc_data_3_16_56_46_sva;
  reg [44:0] buf_acc_data_14_1_45_1_sva;
  reg buf_acc_data_14_1_0_sva;
  reg [10:0] buf_acc_data_14_1_56_46_sva;
  reg [44:0] buf_acc_data_3_15_45_1_sva;
  reg buf_acc_data_3_15_0_sva;
  reg [10:0] buf_acc_data_3_15_56_46_sva;
  reg [44:0] buf_acc_data_14_2_45_1_sva;
  reg buf_acc_data_14_2_0_sva;
  reg [10:0] buf_acc_data_14_2_56_46_sva;
  reg [44:0] buf_acc_data_3_14_45_1_sva;
  reg buf_acc_data_3_14_0_sva;
  reg [10:0] buf_acc_data_3_14_56_46_sva;
  reg [44:0] buf_acc_data_14_3_45_1_sva;
  reg buf_acc_data_14_3_0_sva;
  reg [10:0] buf_acc_data_14_3_56_46_sva;
  reg [44:0] buf_acc_data_3_13_45_1_sva;
  reg buf_acc_data_3_13_0_sva;
  reg [10:0] buf_acc_data_3_13_56_46_sva;
  reg [44:0] buf_acc_data_14_4_45_1_sva;
  reg buf_acc_data_14_4_0_sva;
  reg [10:0] buf_acc_data_14_4_56_46_sva;
  reg [44:0] buf_acc_data_3_12_45_1_sva;
  reg buf_acc_data_3_12_0_sva;
  reg [10:0] buf_acc_data_3_12_56_46_sva;
  reg [44:0] buf_acc_data_14_5_45_1_sva;
  reg buf_acc_data_14_5_0_sva;
  reg [10:0] buf_acc_data_14_5_56_46_sva;
  reg [44:0] buf_acc_data_3_11_45_1_sva;
  reg buf_acc_data_3_11_0_sva;
  reg [10:0] buf_acc_data_3_11_56_46_sva;
  reg [44:0] buf_acc_data_14_6_45_1_sva;
  reg buf_acc_data_14_6_0_sva;
  reg [10:0] buf_acc_data_14_6_56_46_sva;
  reg [44:0] buf_acc_data_3_10_45_1_sva;
  reg buf_acc_data_3_10_0_sva;
  reg [10:0] buf_acc_data_3_10_56_46_sva;
  reg [44:0] buf_acc_data_14_7_45_1_sva;
  reg buf_acc_data_14_7_0_sva;
  reg [10:0] buf_acc_data_14_7_56_46_sva;
  reg [44:0] buf_acc_data_3_9_45_1_sva;
  reg buf_acc_data_3_9_0_sva;
  reg [10:0] buf_acc_data_3_9_56_46_sva;
  reg [44:0] buf_acc_data_14_8_45_1_sva;
  reg buf_acc_data_14_8_0_sva;
  reg [10:0] buf_acc_data_14_8_56_46_sva;
  reg [44:0] buf_acc_data_3_8_45_1_sva;
  reg buf_acc_data_3_8_0_sva;
  reg [10:0] buf_acc_data_3_8_56_46_sva;
  reg [44:0] buf_acc_data_14_9_45_1_sva;
  reg buf_acc_data_14_9_0_sva;
  reg [10:0] buf_acc_data_14_9_56_46_sva;
  reg [44:0] buf_acc_data_3_7_45_1_sva;
  reg buf_acc_data_3_7_0_sva;
  reg [10:0] buf_acc_data_3_7_56_46_sva;
  reg [44:0] buf_acc_data_14_10_45_1_sva;
  reg buf_acc_data_14_10_0_sva;
  reg [10:0] buf_acc_data_14_10_56_46_sva;
  reg [44:0] buf_acc_data_3_6_45_1_sva;
  reg buf_acc_data_3_6_0_sva;
  reg [10:0] buf_acc_data_3_6_56_46_sva;
  reg [44:0] buf_acc_data_14_11_45_1_sva;
  reg buf_acc_data_14_11_0_sva;
  reg [10:0] buf_acc_data_14_11_56_46_sva;
  reg [44:0] buf_acc_data_3_5_45_1_sva;
  reg buf_acc_data_3_5_0_sva;
  reg [10:0] buf_acc_data_3_5_56_46_sva;
  reg [44:0] buf_acc_data_14_12_45_1_sva;
  reg buf_acc_data_14_12_0_sva;
  reg [10:0] buf_acc_data_14_12_56_46_sva;
  reg [44:0] buf_acc_data_3_4_45_1_sva;
  reg buf_acc_data_3_4_0_sva;
  reg [10:0] buf_acc_data_3_4_56_46_sva;
  reg [44:0] buf_acc_data_14_13_45_1_sva;
  reg buf_acc_data_14_13_0_sva;
  reg [10:0] buf_acc_data_14_13_56_46_sva;
  reg [44:0] buf_acc_data_3_3_45_1_sva;
  reg buf_acc_data_3_3_0_sva;
  reg [10:0] buf_acc_data_3_3_56_46_sva;
  reg [44:0] buf_acc_data_14_14_45_1_sva;
  reg buf_acc_data_14_14_0_sva;
  reg [10:0] buf_acc_data_14_14_56_46_sva;
  reg [44:0] buf_acc_data_3_2_45_1_sva;
  reg buf_acc_data_3_2_0_sva;
  reg [10:0] buf_acc_data_3_2_56_46_sva;
  reg [44:0] buf_acc_data_14_15_45_1_sva;
  reg buf_acc_data_14_15_0_sva;
  reg [10:0] buf_acc_data_14_15_56_46_sva;
  reg [44:0] buf_acc_data_3_1_45_1_sva;
  reg buf_acc_data_3_1_0_sva;
  reg [10:0] buf_acc_data_3_1_56_46_sva;
  reg [44:0] buf_acc_data_14_16_45_1_sva;
  reg buf_acc_data_14_16_0_sva;
  reg [10:0] buf_acc_data_14_16_56_46_sva;
  reg [44:0] buf_acc_data_3_0_45_1_sva;
  reg buf_acc_data_3_0_0_sva;
  reg [10:0] buf_acc_data_3_0_56_46_sva;
  reg [44:0] buf_acc_data_14_17_45_1_sva;
  reg buf_acc_data_14_17_0_sva;
  reg [10:0] buf_acc_data_14_17_56_46_sva;
  reg [44:0] buf_acc_data_2_17_45_1_sva;
  reg buf_acc_data_2_17_0_sva;
  reg [10:0] buf_acc_data_2_17_56_46_sva;
  reg [44:0] buf_acc_data_15_0_45_1_sva;
  reg buf_acc_data_15_0_0_sva;
  reg [10:0] buf_acc_data_15_0_56_46_sva;
  reg [44:0] buf_acc_data_2_16_45_1_sva;
  reg buf_acc_data_2_16_0_sva;
  reg [10:0] buf_acc_data_2_16_56_46_sva;
  reg [44:0] buf_acc_data_15_1_45_1_sva;
  reg buf_acc_data_15_1_0_sva;
  reg [10:0] buf_acc_data_15_1_56_46_sva;
  reg [44:0] buf_acc_data_2_15_45_1_sva;
  reg buf_acc_data_2_15_0_sva;
  reg [10:0] buf_acc_data_2_15_56_46_sva;
  reg [44:0] buf_acc_data_15_2_45_1_sva;
  reg buf_acc_data_15_2_0_sva;
  reg [10:0] buf_acc_data_15_2_56_46_sva;
  reg [44:0] buf_acc_data_2_14_45_1_sva;
  reg buf_acc_data_2_14_0_sva;
  reg [10:0] buf_acc_data_2_14_56_46_sva;
  reg [44:0] buf_acc_data_15_3_45_1_sva;
  reg buf_acc_data_15_3_0_sva;
  reg [10:0] buf_acc_data_15_3_56_46_sva;
  reg [44:0] buf_acc_data_2_13_45_1_sva;
  reg buf_acc_data_2_13_0_sva;
  reg [10:0] buf_acc_data_2_13_56_46_sva;
  reg [44:0] buf_acc_data_15_4_45_1_sva;
  reg buf_acc_data_15_4_0_sva;
  reg [10:0] buf_acc_data_15_4_56_46_sva;
  reg [44:0] buf_acc_data_2_12_45_1_sva;
  reg buf_acc_data_2_12_0_sva;
  reg [10:0] buf_acc_data_2_12_56_46_sva;
  reg [44:0] buf_acc_data_15_5_45_1_sva;
  reg buf_acc_data_15_5_0_sva;
  reg [10:0] buf_acc_data_15_5_56_46_sva;
  reg [44:0] buf_acc_data_2_11_45_1_sva;
  reg buf_acc_data_2_11_0_sva;
  reg [10:0] buf_acc_data_2_11_56_46_sva;
  reg [44:0] buf_acc_data_15_6_45_1_sva;
  reg buf_acc_data_15_6_0_sva;
  reg [10:0] buf_acc_data_15_6_56_46_sva;
  reg [44:0] buf_acc_data_2_10_45_1_sva;
  reg buf_acc_data_2_10_0_sva;
  reg [10:0] buf_acc_data_2_10_56_46_sva;
  reg [44:0] buf_acc_data_15_7_45_1_sva;
  reg buf_acc_data_15_7_0_sva;
  reg [10:0] buf_acc_data_15_7_56_46_sva;
  reg [44:0] buf_acc_data_2_9_45_1_sva;
  reg buf_acc_data_2_9_0_sva;
  reg [10:0] buf_acc_data_2_9_56_46_sva;
  reg [44:0] buf_acc_data_15_8_45_1_sva;
  reg buf_acc_data_15_8_0_sva;
  reg [10:0] buf_acc_data_15_8_56_46_sva;
  reg [44:0] buf_acc_data_2_8_45_1_sva;
  reg buf_acc_data_2_8_0_sva;
  reg [10:0] buf_acc_data_2_8_56_46_sva;
  reg [44:0] buf_acc_data_15_9_45_1_sva;
  reg buf_acc_data_15_9_0_sva;
  reg [10:0] buf_acc_data_15_9_56_46_sva;
  reg [44:0] buf_acc_data_2_7_45_1_sva;
  reg buf_acc_data_2_7_0_sva;
  reg [10:0] buf_acc_data_2_7_56_46_sva;
  reg [44:0] buf_acc_data_15_10_45_1_sva;
  reg buf_acc_data_15_10_0_sva;
  reg [10:0] buf_acc_data_15_10_56_46_sva;
  reg [44:0] buf_acc_data_2_6_45_1_sva;
  reg buf_acc_data_2_6_0_sva;
  reg [10:0] buf_acc_data_2_6_56_46_sva;
  reg [44:0] buf_acc_data_15_11_45_1_sva;
  reg buf_acc_data_15_11_0_sva;
  reg [10:0] buf_acc_data_15_11_56_46_sva;
  reg [44:0] buf_acc_data_2_5_45_1_sva;
  reg buf_acc_data_2_5_0_sva;
  reg [10:0] buf_acc_data_2_5_56_46_sva;
  reg [44:0] buf_acc_data_15_12_45_1_sva;
  reg buf_acc_data_15_12_0_sva;
  reg [10:0] buf_acc_data_15_12_56_46_sva;
  reg [44:0] buf_acc_data_2_4_45_1_sva;
  reg buf_acc_data_2_4_0_sva;
  reg [10:0] buf_acc_data_2_4_56_46_sva;
  reg [44:0] buf_acc_data_15_13_45_1_sva;
  reg buf_acc_data_15_13_0_sva;
  reg [10:0] buf_acc_data_15_13_56_46_sva;
  reg [44:0] buf_acc_data_2_3_45_1_sva;
  reg buf_acc_data_2_3_0_sva;
  reg [10:0] buf_acc_data_2_3_56_46_sva;
  reg [44:0] buf_acc_data_15_14_45_1_sva;
  reg buf_acc_data_15_14_0_sva;
  reg [10:0] buf_acc_data_15_14_56_46_sva;
  reg [44:0] buf_acc_data_2_2_45_1_sva;
  reg buf_acc_data_2_2_0_sva;
  reg [10:0] buf_acc_data_2_2_56_46_sva;
  reg [44:0] buf_acc_data_15_15_45_1_sva;
  reg buf_acc_data_15_15_0_sva;
  reg [10:0] buf_acc_data_15_15_56_46_sva;
  reg [44:0] buf_acc_data_2_1_45_1_sva;
  reg buf_acc_data_2_1_0_sva;
  reg [10:0] buf_acc_data_2_1_56_46_sva;
  reg [44:0] buf_acc_data_15_16_45_1_sva;
  reg buf_acc_data_15_16_0_sva;
  reg [10:0] buf_acc_data_15_16_56_46_sva;
  reg [44:0] buf_acc_data_2_0_45_1_sva;
  reg buf_acc_data_2_0_0_sva;
  reg [10:0] buf_acc_data_2_0_56_46_sva;
  reg [44:0] buf_acc_data_15_17_45_1_sva;
  reg buf_acc_data_15_17_0_sva;
  reg [10:0] buf_acc_data_15_17_56_46_sva;
  reg [44:0] buf_acc_data_1_17_45_1_sva;
  reg buf_acc_data_1_17_0_sva;
  reg [10:0] buf_acc_data_1_17_56_46_sva;
  reg [44:0] buf_acc_data_16_0_45_1_sva;
  reg buf_acc_data_16_0_0_sva;
  reg [10:0] buf_acc_data_16_0_56_46_sva;
  reg [44:0] buf_acc_data_1_16_45_1_sva;
  reg buf_acc_data_1_16_0_sva;
  reg [10:0] buf_acc_data_1_16_56_46_sva;
  reg [44:0] buf_acc_data_16_1_45_1_sva;
  reg buf_acc_data_16_1_0_sva;
  reg [10:0] buf_acc_data_16_1_56_46_sva;
  reg [44:0] buf_acc_data_1_15_45_1_sva;
  reg buf_acc_data_1_15_0_sva;
  reg [10:0] buf_acc_data_1_15_56_46_sva;
  reg [44:0] buf_acc_data_16_2_45_1_sva;
  reg buf_acc_data_16_2_0_sva;
  reg [10:0] buf_acc_data_16_2_56_46_sva;
  reg [44:0] buf_acc_data_1_14_45_1_sva;
  reg buf_acc_data_1_14_0_sva;
  reg [10:0] buf_acc_data_1_14_56_46_sva;
  reg [44:0] buf_acc_data_16_3_45_1_sva;
  reg buf_acc_data_16_3_0_sva;
  reg [10:0] buf_acc_data_16_3_56_46_sva;
  reg [44:0] buf_acc_data_1_13_45_1_sva;
  reg buf_acc_data_1_13_0_sva;
  reg [10:0] buf_acc_data_1_13_56_46_sva;
  reg [44:0] buf_acc_data_16_4_45_1_sva;
  reg buf_acc_data_16_4_0_sva;
  reg [10:0] buf_acc_data_16_4_56_46_sva;
  reg [44:0] buf_acc_data_1_12_45_1_sva;
  reg buf_acc_data_1_12_0_sva;
  reg [10:0] buf_acc_data_1_12_56_46_sva;
  reg [44:0] buf_acc_data_16_5_45_1_sva;
  reg buf_acc_data_16_5_0_sva;
  reg [10:0] buf_acc_data_16_5_56_46_sva;
  reg [44:0] buf_acc_data_1_11_45_1_sva;
  reg buf_acc_data_1_11_0_sva;
  reg [10:0] buf_acc_data_1_11_56_46_sva;
  reg [44:0] buf_acc_data_16_6_45_1_sva;
  reg buf_acc_data_16_6_0_sva;
  reg [10:0] buf_acc_data_16_6_56_46_sva;
  reg [44:0] buf_acc_data_1_10_45_1_sva;
  reg buf_acc_data_1_10_0_sva;
  reg [10:0] buf_acc_data_1_10_56_46_sva;
  reg [44:0] buf_acc_data_16_7_45_1_sva;
  reg buf_acc_data_16_7_0_sva;
  reg [10:0] buf_acc_data_16_7_56_46_sva;
  reg [44:0] buf_acc_data_1_9_45_1_sva;
  reg buf_acc_data_1_9_0_sva;
  reg [10:0] buf_acc_data_1_9_56_46_sva;
  reg [44:0] buf_acc_data_16_8_45_1_sva;
  reg buf_acc_data_16_8_0_sva;
  reg [10:0] buf_acc_data_16_8_56_46_sva;
  reg [44:0] buf_acc_data_1_8_45_1_sva;
  reg buf_acc_data_1_8_0_sva;
  reg [10:0] buf_acc_data_1_8_56_46_sva;
  reg [44:0] buf_acc_data_16_9_45_1_sva;
  reg buf_acc_data_16_9_0_sva;
  reg [10:0] buf_acc_data_16_9_56_46_sva;
  reg [44:0] buf_acc_data_1_7_45_1_sva;
  reg buf_acc_data_1_7_0_sva;
  reg [10:0] buf_acc_data_1_7_56_46_sva;
  reg [44:0] buf_acc_data_16_10_45_1_sva;
  reg buf_acc_data_16_10_0_sva;
  reg [10:0] buf_acc_data_16_10_56_46_sva;
  reg [44:0] buf_acc_data_1_6_45_1_sva;
  reg buf_acc_data_1_6_0_sva;
  reg [10:0] buf_acc_data_1_6_56_46_sva;
  reg [44:0] buf_acc_data_16_11_45_1_sva;
  reg buf_acc_data_16_11_0_sva;
  reg [10:0] buf_acc_data_16_11_56_46_sva;
  reg [44:0] buf_acc_data_1_5_45_1_sva;
  reg buf_acc_data_1_5_0_sva;
  reg [10:0] buf_acc_data_1_5_56_46_sva;
  reg [44:0] buf_acc_data_16_12_45_1_sva;
  reg buf_acc_data_16_12_0_sva;
  reg [10:0] buf_acc_data_16_12_56_46_sva;
  reg [44:0] buf_acc_data_1_4_45_1_sva;
  reg buf_acc_data_1_4_0_sva;
  reg [10:0] buf_acc_data_1_4_56_46_sva;
  reg [44:0] buf_acc_data_16_13_45_1_sva;
  reg buf_acc_data_16_13_0_sva;
  reg [10:0] buf_acc_data_16_13_56_46_sva;
  reg [44:0] buf_acc_data_1_3_45_1_sva;
  reg buf_acc_data_1_3_0_sva;
  reg [10:0] buf_acc_data_1_3_56_46_sva;
  reg [44:0] buf_acc_data_16_14_45_1_sva;
  reg buf_acc_data_16_14_0_sva;
  reg [10:0] buf_acc_data_16_14_56_46_sva;
  reg [44:0] buf_acc_data_1_2_45_1_sva;
  reg buf_acc_data_1_2_0_sva;
  reg [10:0] buf_acc_data_1_2_56_46_sva;
  reg [44:0] buf_acc_data_16_15_45_1_sva;
  reg buf_acc_data_16_15_0_sva;
  reg [10:0] buf_acc_data_16_15_56_46_sva;
  reg [44:0] buf_acc_data_1_1_45_1_sva;
  reg buf_acc_data_1_1_0_sva;
  reg [10:0] buf_acc_data_1_1_56_46_sva;
  reg [44:0] buf_acc_data_16_16_45_1_sva;
  reg buf_acc_data_16_16_0_sva;
  reg [10:0] buf_acc_data_16_16_56_46_sva;
  reg [44:0] buf_acc_data_1_0_45_1_sva;
  reg buf_acc_data_1_0_0_sva;
  reg [10:0] buf_acc_data_1_0_56_46_sva;
  reg [44:0] buf_acc_data_16_17_45_1_sva;
  reg buf_acc_data_16_17_0_sva;
  reg [10:0] buf_acc_data_16_17_56_46_sva;
  reg [44:0] buf_acc_data_0_17_45_1_sva;
  reg buf_acc_data_0_17_0_sva;
  reg [10:0] buf_acc_data_0_17_56_46_sva;
  reg [44:0] buf_acc_data_17_0_45_1_sva;
  reg buf_acc_data_17_0_0_sva;
  reg [10:0] buf_acc_data_17_0_56_46_sva;
  reg [44:0] buf_acc_data_0_16_45_1_sva;
  reg buf_acc_data_0_16_0_sva;
  reg [10:0] buf_acc_data_0_16_56_46_sva;
  reg [44:0] buf_acc_data_17_1_45_1_sva;
  reg buf_acc_data_17_1_0_sva;
  reg [10:0] buf_acc_data_17_1_56_46_sva;
  reg [44:0] buf_acc_data_0_15_45_1_sva;
  reg buf_acc_data_0_15_0_sva;
  reg [10:0] buf_acc_data_0_15_56_46_sva;
  reg [44:0] buf_acc_data_17_2_45_1_sva;
  reg buf_acc_data_17_2_0_sva;
  reg [10:0] buf_acc_data_17_2_56_46_sva;
  reg [44:0] buf_acc_data_0_14_45_1_sva;
  reg buf_acc_data_0_14_0_sva;
  reg [10:0] buf_acc_data_0_14_56_46_sva;
  reg [44:0] buf_acc_data_17_3_45_1_sva;
  reg buf_acc_data_17_3_0_sva;
  reg [10:0] buf_acc_data_17_3_56_46_sva;
  reg [44:0] buf_acc_data_0_13_45_1_sva;
  reg buf_acc_data_0_13_0_sva;
  reg [10:0] buf_acc_data_0_13_56_46_sva;
  reg [44:0] buf_acc_data_17_4_45_1_sva;
  reg buf_acc_data_17_4_0_sva;
  reg [10:0] buf_acc_data_17_4_56_46_sva;
  reg [44:0] buf_acc_data_0_12_45_1_sva;
  reg buf_acc_data_0_12_0_sva;
  reg [10:0] buf_acc_data_0_12_56_46_sva;
  reg [44:0] buf_acc_data_17_5_45_1_sva;
  reg buf_acc_data_17_5_0_sva;
  reg [10:0] buf_acc_data_17_5_56_46_sva;
  reg [44:0] buf_acc_data_0_11_45_1_sva;
  reg buf_acc_data_0_11_0_sva;
  reg [10:0] buf_acc_data_0_11_56_46_sva;
  reg [44:0] buf_acc_data_17_6_45_1_sva;
  reg buf_acc_data_17_6_0_sva;
  reg [10:0] buf_acc_data_17_6_56_46_sva;
  reg [44:0] buf_acc_data_0_10_45_1_sva;
  reg buf_acc_data_0_10_0_sva;
  reg [10:0] buf_acc_data_0_10_56_46_sva;
  reg [44:0] buf_acc_data_17_7_45_1_sva;
  reg buf_acc_data_17_7_0_sva;
  reg [10:0] buf_acc_data_17_7_56_46_sva;
  reg [44:0] buf_acc_data_0_9_45_1_sva;
  reg buf_acc_data_0_9_0_sva;
  reg [10:0] buf_acc_data_0_9_56_46_sva;
  reg [44:0] buf_acc_data_17_8_45_1_sva;
  reg buf_acc_data_17_8_0_sva;
  reg [10:0] buf_acc_data_17_8_56_46_sva;
  reg [44:0] buf_acc_data_0_8_45_1_sva;
  reg buf_acc_data_0_8_0_sva;
  reg [10:0] buf_acc_data_0_8_56_46_sva;
  reg [44:0] buf_acc_data_17_9_45_1_sva;
  reg buf_acc_data_17_9_0_sva;
  reg [10:0] buf_acc_data_17_9_56_46_sva;
  reg [44:0] buf_acc_data_0_7_45_1_sva;
  reg buf_acc_data_0_7_0_sva;
  reg [10:0] buf_acc_data_0_7_56_46_sva;
  reg [44:0] buf_acc_data_17_10_45_1_sva;
  reg buf_acc_data_17_10_0_sva;
  reg [10:0] buf_acc_data_17_10_56_46_sva;
  reg [44:0] buf_acc_data_0_6_45_1_sva;
  reg buf_acc_data_0_6_0_sva;
  reg [10:0] buf_acc_data_0_6_56_46_sva;
  reg [44:0] buf_acc_data_17_11_45_1_sva;
  reg buf_acc_data_17_11_0_sva;
  reg [10:0] buf_acc_data_17_11_56_46_sva;
  reg [44:0] buf_acc_data_0_5_45_1_sva;
  reg buf_acc_data_0_5_0_sva;
  reg [10:0] buf_acc_data_0_5_56_46_sva;
  reg [44:0] buf_acc_data_17_12_45_1_sva;
  reg buf_acc_data_17_12_0_sva;
  reg [10:0] buf_acc_data_17_12_56_46_sva;
  reg [44:0] buf_acc_data_0_4_45_1_sva;
  reg buf_acc_data_0_4_0_sva;
  reg [10:0] buf_acc_data_0_4_56_46_sva;
  reg [44:0] buf_acc_data_17_13_45_1_sva;
  reg buf_acc_data_17_13_0_sva;
  reg [10:0] buf_acc_data_17_13_56_46_sva;
  reg [44:0] buf_acc_data_0_3_45_1_sva;
  reg buf_acc_data_0_3_0_sva;
  reg [10:0] buf_acc_data_0_3_56_46_sva;
  reg [44:0] buf_acc_data_17_14_45_1_sva;
  reg buf_acc_data_17_14_0_sva;
  reg [10:0] buf_acc_data_17_14_56_46_sva;
  reg [44:0] buf_acc_data_0_2_45_1_sva;
  reg buf_acc_data_0_2_0_sva;
  reg [10:0] buf_acc_data_0_2_56_46_sva;
  reg [44:0] buf_acc_data_17_15_45_1_sva;
  reg buf_acc_data_17_15_0_sva;
  reg [10:0] buf_acc_data_17_15_56_46_sva;
  reg [44:0] buf_acc_data_0_1_45_1_sva;
  reg buf_acc_data_0_1_0_sva;
  reg [10:0] buf_acc_data_0_1_56_46_sva;
  reg [44:0] buf_acc_data_17_16_45_1_sva;
  reg buf_acc_data_17_16_0_sva;
  reg [10:0] buf_acc_data_17_16_56_46_sva;
  reg [44:0] buf_acc_data_0_0_45_1_sva;
  reg buf_acc_data_0_0_0_sva;
  reg [10:0] buf_acc_data_0_0_56_46_sva;
  reg [44:0] buf_acc_data_17_17_45_1_sva;
  reg buf_acc_data_17_17_0_sva;
  reg [10:0] buf_acc_data_17_17_56_46_sva;
  reg [7:0] pad_sva;
  reg [6:0] n_w_in_acc_psp_sva;
  wire [7:0] nl_n_w_in_acc_psp_sva;
  reg [6:0] n_h_in_acc_psp_sva;
  wire [7:0] nl_n_h_in_acc_psp_sva;
  reg [7:0] n_w_out_lpi_1_dfm;
  reg [7:0] n_h_out_lpi_1_dfm;
  reg [15:0] dma_read_data_length_mul_4_cse_sva;
  reg [15:0] dma_read_data_length_sva;
  reg [15:0] dma_write_data_length_sva;
  wire [23:0] nl_dma_write_data_length_sva;
  reg [15:0] dma_read_info_index_15_0_lpi_2_dfm;
  reg [15:0] LOAD_LOOP_i_lpi_2_dfm_2;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_2;
  reg CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_dfm_1;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_dfm_1;
  reg CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_dfm_1;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1;
  reg [4:0] PADDING_LOOP_for_row_4_0_lpi_2_dfm_5;
  reg [4:0] PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4;
  reg [4:0] CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4;
  reg [13:0] STORE_LOOP_i_13_0_lpi_2_dfm_2;
  reg lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3;
  reg lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_1;
  reg lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1;
  reg lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1;
  reg lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1;
  reg BATCH_LOOP_stage_v_1;
  reg PADDING_LOOP_for_for_land_2_lpi_2_dfm_st;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st;
  reg [10:0] CONVOLUTION_LOOP_for_for_for_else_mux_itm;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_else_mux_972_itm;
  reg CONVOLUTION_LOOP_for_for_for_else_mux_973_itm;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm;
  reg exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st;
  reg exit_CONVOLUTION_LOOP_lpi_2_dfm_2_1;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1;
  reg [15:0] LOAD_LOOP_i_sva_1_1;
  reg PADDING_LOOP_for_for_land_2_lpi_2_dfm_1;
  reg [13:0] PADDING_LOOP_for_for_index_in_acc_itm_1;
  wire [14:0] nl_PADDING_LOOP_for_for_index_in_acc_itm_1;
  reg [15:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1;
  wire [16:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1;
  reg [13:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1;
  wire [14:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_1;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_1;
  reg [13:0] CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1;
  wire [14:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1;
  reg [13:0] CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2;
  reg [13:0] STORE_LOOP_data_asn_itm_1;
  reg STORE_LOOP_and_30_itm_1;
  reg STORE_LOOP_and_32_itm_1;
  reg [4:0] CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0;
  reg [231:0] conf_info_crt_sva_231_0;
  reg [3:0] BATCH_LOOP_b_4_0_sva_3_0;
  reg [4:0] PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0;
  reg [4:0] CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0;
  reg [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0;
  reg CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_1_0;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_7_3;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_2_0;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_7_3;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_0;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_8_2;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_8_1;
  reg lfst_exit_STORE_LOOP_lpi_2_dfm_8_0;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_7_3;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_2_0;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0;
  wire [4:0] PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0_mx1w0;
  wire [4:0] CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0_mx1w0;
  wire PADDING_LOOP_for_for_land_2_lpi_2_dfm_mx1w0;
  wire PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1_mx0c1;
  wire exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1_mx0c1;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1_mx0c1;
  wire exit_BATCH_LOOP_lpi_2_dfm_2_mx1w0;
  wire [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0_mx1w0;
  wire CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1;
  wire [44:0] CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_mx1;
  wire CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_mx0w0;
  wire [44:0] CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_mx0w0;
  wire [10:0] CONVOLUTION_LOOP_for_for_for_else_mux_itm_mx0w0;
  wire exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0;
  wire [15:0] LOAD_LOOP_i_lpi_2_dfm_2_mx0w0;
  wire [4:0] PADDING_LOOP_for_row_4_0_lpi_2_dfm_5_mx0w0;
  wire lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0;
  wire [4:0] PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4_mx0w0;
  wire lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0;
  wire [4:0] CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5_mx0w0;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5_mx0w0;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2_mx0w0;
  wire CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1_mx0c1;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3_mx0w0;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4_mx0w0;
  wire [13:0] STORE_LOOP_i_13_0_lpi_2_dfm_2_mx0w0;
  wire [7:0] if_acc_4_cse_1;
  wire [8:0] nl_if_acc_4_cse_1;
  wire [10:0] else_acc_2_psp_sva_1;
  wire [11:0] nl_else_acc_2_psp_sva_1;
  wire [10:0] else_acc_psp_sva_1;
  wire [11:0] nl_else_acc_psp_sva_1;
  wire BATCH_LOOP_stage_v_2_mx0c0;
  wire BATCH_LOOP_stage_v_3_mx0c0;
  wire LOAD_LOOP_i_lpi_2_mx0c1;
  wire [7:0] asn_3_mx0w1;
  wire [8:0] nl_asn_3_mx0w1;
  wire [7:0] asn_1_mx0w0;
  wire [8:0] nl_asn_1_mx0w0;
  wire [7:0] asn_mx0w1;
  wire [8:0] nl_asn_mx0w1;
  wire buf_acc_data_17_17_0_sva_mx0;
  wire [44:0] buf_acc_data_17_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_17_56_46_sva_mx0;
  wire buf_acc_data_0_0_0_sva_mx0;
  wire [44:0] buf_acc_data_0_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_0_56_46_sva_mx0;
  wire buf_acc_data_17_16_0_sva_mx0;
  wire [44:0] buf_acc_data_17_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_16_56_46_sva_mx0;
  wire buf_acc_data_0_1_0_sva_mx0;
  wire [44:0] buf_acc_data_0_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_1_56_46_sva_mx0;
  wire buf_acc_data_17_15_0_sva_mx0;
  wire [44:0] buf_acc_data_17_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_15_56_46_sva_mx0;
  wire buf_acc_data_0_2_0_sva_mx0;
  wire [44:0] buf_acc_data_0_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_2_56_46_sva_mx0;
  wire buf_acc_data_17_14_0_sva_mx0;
  wire [44:0] buf_acc_data_17_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_14_56_46_sva_mx0;
  wire buf_acc_data_0_3_0_sva_mx0;
  wire [44:0] buf_acc_data_0_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_3_56_46_sva_mx0;
  wire buf_acc_data_17_13_0_sva_mx0;
  wire [44:0] buf_acc_data_17_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_13_56_46_sva_mx0;
  wire buf_acc_data_0_4_0_sva_mx0;
  wire [44:0] buf_acc_data_0_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_4_56_46_sva_mx0;
  wire buf_acc_data_17_12_0_sva_mx0;
  wire [44:0] buf_acc_data_17_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_12_56_46_sva_mx0;
  wire buf_acc_data_0_5_0_sva_mx0;
  wire [44:0] buf_acc_data_0_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_5_56_46_sva_mx0;
  wire buf_acc_data_17_11_0_sva_mx0;
  wire [44:0] buf_acc_data_17_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_11_56_46_sva_mx0;
  wire buf_acc_data_0_6_0_sva_mx0;
  wire [44:0] buf_acc_data_0_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_6_56_46_sva_mx0;
  wire buf_acc_data_17_10_0_sva_mx0;
  wire [44:0] buf_acc_data_17_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_10_56_46_sva_mx0;
  wire buf_acc_data_0_7_0_sva_mx0;
  wire [44:0] buf_acc_data_0_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_7_56_46_sva_mx0;
  wire buf_acc_data_17_9_0_sva_mx0;
  wire [44:0] buf_acc_data_17_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_9_56_46_sva_mx0;
  wire buf_acc_data_0_8_0_sva_mx0;
  wire [44:0] buf_acc_data_0_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_8_56_46_sva_mx0;
  wire buf_acc_data_17_8_0_sva_mx0;
  wire [44:0] buf_acc_data_17_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_8_56_46_sva_mx0;
  wire buf_acc_data_0_9_0_sva_mx0;
  wire [44:0] buf_acc_data_0_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_9_56_46_sva_mx0;
  wire buf_acc_data_17_7_0_sva_mx0;
  wire [44:0] buf_acc_data_17_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_7_56_46_sva_mx0;
  wire buf_acc_data_0_10_0_sva_mx0;
  wire [44:0] buf_acc_data_0_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_10_56_46_sva_mx0;
  wire buf_acc_data_17_6_0_sva_mx0;
  wire [44:0] buf_acc_data_17_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_6_56_46_sva_mx0;
  wire buf_acc_data_0_11_0_sva_mx0;
  wire [44:0] buf_acc_data_0_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_11_56_46_sva_mx0;
  wire buf_acc_data_17_5_0_sva_mx0;
  wire [44:0] buf_acc_data_17_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_5_56_46_sva_mx0;
  wire buf_acc_data_0_12_0_sva_mx0;
  wire [44:0] buf_acc_data_0_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_12_56_46_sva_mx0;
  wire buf_acc_data_17_4_0_sva_mx0;
  wire [44:0] buf_acc_data_17_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_4_56_46_sva_mx0;
  wire buf_acc_data_0_13_0_sva_mx0;
  wire [44:0] buf_acc_data_0_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_13_56_46_sva_mx0;
  wire buf_acc_data_17_3_0_sva_mx0;
  wire [44:0] buf_acc_data_17_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_3_56_46_sva_mx0;
  wire buf_acc_data_0_14_0_sva_mx0;
  wire [44:0] buf_acc_data_0_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_14_56_46_sva_mx0;
  wire buf_acc_data_17_2_0_sva_mx0;
  wire [44:0] buf_acc_data_17_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_2_56_46_sva_mx0;
  wire buf_acc_data_0_15_0_sva_mx0;
  wire [44:0] buf_acc_data_0_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_15_56_46_sva_mx0;
  wire buf_acc_data_17_1_0_sva_mx0;
  wire [44:0] buf_acc_data_17_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_1_56_46_sva_mx0;
  wire buf_acc_data_0_16_0_sva_mx0;
  wire [44:0] buf_acc_data_0_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_16_56_46_sva_mx0;
  wire buf_acc_data_17_0_0_sva_mx0;
  wire [44:0] buf_acc_data_17_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_17_0_56_46_sva_mx0;
  wire buf_acc_data_0_17_0_sva_mx0;
  wire [44:0] buf_acc_data_0_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_0_17_56_46_sva_mx0;
  wire buf_acc_data_16_17_0_sva_mx0;
  wire [44:0] buf_acc_data_16_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_17_56_46_sva_mx0;
  wire buf_acc_data_1_0_0_sva_mx0;
  wire [44:0] buf_acc_data_1_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_0_56_46_sva_mx0;
  wire buf_acc_data_16_16_0_sva_mx0;
  wire [44:0] buf_acc_data_16_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_16_56_46_sva_mx0;
  wire buf_acc_data_1_1_0_sva_mx0;
  wire [44:0] buf_acc_data_1_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_1_56_46_sva_mx0;
  wire buf_acc_data_16_15_0_sva_mx0;
  wire [44:0] buf_acc_data_16_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_15_56_46_sva_mx0;
  wire buf_acc_data_1_2_0_sva_mx0;
  wire [44:0] buf_acc_data_1_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_2_56_46_sva_mx0;
  wire buf_acc_data_16_14_0_sva_mx0;
  wire [44:0] buf_acc_data_16_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_14_56_46_sva_mx0;
  wire buf_acc_data_1_3_0_sva_mx0;
  wire [44:0] buf_acc_data_1_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_3_56_46_sva_mx0;
  wire buf_acc_data_16_13_0_sva_mx0;
  wire [44:0] buf_acc_data_16_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_13_56_46_sva_mx0;
  wire buf_acc_data_1_4_0_sva_mx0;
  wire [44:0] buf_acc_data_1_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_4_56_46_sva_mx0;
  wire buf_acc_data_16_12_0_sva_mx0;
  wire [44:0] buf_acc_data_16_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_12_56_46_sva_mx0;
  wire buf_acc_data_1_5_0_sva_mx0;
  wire [44:0] buf_acc_data_1_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_5_56_46_sva_mx0;
  wire buf_acc_data_16_11_0_sva_mx0;
  wire [44:0] buf_acc_data_16_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_11_56_46_sva_mx0;
  wire buf_acc_data_1_6_0_sva_mx0;
  wire [44:0] buf_acc_data_1_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_6_56_46_sva_mx0;
  wire buf_acc_data_16_10_0_sva_mx0;
  wire [44:0] buf_acc_data_16_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_10_56_46_sva_mx0;
  wire buf_acc_data_1_7_0_sva_mx0;
  wire [44:0] buf_acc_data_1_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_7_56_46_sva_mx0;
  wire buf_acc_data_16_9_0_sva_mx0;
  wire [44:0] buf_acc_data_16_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_9_56_46_sva_mx0;
  wire buf_acc_data_1_8_0_sva_mx0;
  wire [44:0] buf_acc_data_1_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_8_56_46_sva_mx0;
  wire buf_acc_data_16_8_0_sva_mx0;
  wire [44:0] buf_acc_data_16_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_8_56_46_sva_mx0;
  wire buf_acc_data_1_9_0_sva_mx0;
  wire [44:0] buf_acc_data_1_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_9_56_46_sva_mx0;
  wire buf_acc_data_16_7_0_sva_mx0;
  wire [44:0] buf_acc_data_16_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_7_56_46_sva_mx0;
  wire buf_acc_data_1_10_0_sva_mx0;
  wire [44:0] buf_acc_data_1_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_10_56_46_sva_mx0;
  wire buf_acc_data_16_6_0_sva_mx0;
  wire [44:0] buf_acc_data_16_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_6_56_46_sva_mx0;
  wire buf_acc_data_1_11_0_sva_mx0;
  wire [44:0] buf_acc_data_1_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_11_56_46_sva_mx0;
  wire buf_acc_data_16_5_0_sva_mx0;
  wire [44:0] buf_acc_data_16_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_5_56_46_sva_mx0;
  wire buf_acc_data_1_12_0_sva_mx0;
  wire [44:0] buf_acc_data_1_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_12_56_46_sva_mx0;
  wire buf_acc_data_16_4_0_sva_mx0;
  wire [44:0] buf_acc_data_16_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_4_56_46_sva_mx0;
  wire buf_acc_data_1_13_0_sva_mx0;
  wire [44:0] buf_acc_data_1_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_13_56_46_sva_mx0;
  wire buf_acc_data_16_3_0_sva_mx0;
  wire [44:0] buf_acc_data_16_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_3_56_46_sva_mx0;
  wire buf_acc_data_1_14_0_sva_mx0;
  wire [44:0] buf_acc_data_1_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_14_56_46_sva_mx0;
  wire buf_acc_data_16_2_0_sva_mx0;
  wire [44:0] buf_acc_data_16_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_2_56_46_sva_mx0;
  wire buf_acc_data_1_15_0_sva_mx0;
  wire [44:0] buf_acc_data_1_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_15_56_46_sva_mx0;
  wire buf_acc_data_16_1_0_sva_mx0;
  wire [44:0] buf_acc_data_16_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_1_56_46_sva_mx0;
  wire buf_acc_data_1_16_0_sva_mx0;
  wire [44:0] buf_acc_data_1_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_16_56_46_sva_mx0;
  wire buf_acc_data_16_0_0_sva_mx0;
  wire [44:0] buf_acc_data_16_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_16_0_56_46_sva_mx0;
  wire buf_acc_data_1_17_0_sva_mx0;
  wire [44:0] buf_acc_data_1_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_1_17_56_46_sva_mx0;
  wire buf_acc_data_15_17_0_sva_mx0;
  wire [44:0] buf_acc_data_15_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_17_56_46_sva_mx0;
  wire buf_acc_data_2_0_0_sva_mx0;
  wire [44:0] buf_acc_data_2_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_0_56_46_sva_mx0;
  wire buf_acc_data_15_16_0_sva_mx0;
  wire [44:0] buf_acc_data_15_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_16_56_46_sva_mx0;
  wire buf_acc_data_2_1_0_sva_mx0;
  wire [44:0] buf_acc_data_2_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_1_56_46_sva_mx0;
  wire buf_acc_data_15_15_0_sva_mx0;
  wire [44:0] buf_acc_data_15_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_15_56_46_sva_mx0;
  wire buf_acc_data_2_2_0_sva_mx0;
  wire [44:0] buf_acc_data_2_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_2_56_46_sva_mx0;
  wire buf_acc_data_15_14_0_sva_mx0;
  wire [44:0] buf_acc_data_15_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_14_56_46_sva_mx0;
  wire buf_acc_data_2_3_0_sva_mx0;
  wire [44:0] buf_acc_data_2_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_3_56_46_sva_mx0;
  wire buf_acc_data_15_13_0_sva_mx0;
  wire [44:0] buf_acc_data_15_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_13_56_46_sva_mx0;
  wire buf_acc_data_2_4_0_sva_mx0;
  wire [44:0] buf_acc_data_2_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_4_56_46_sva_mx0;
  wire buf_acc_data_15_12_0_sva_mx0;
  wire [44:0] buf_acc_data_15_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_12_56_46_sva_mx0;
  wire buf_acc_data_2_5_0_sva_mx0;
  wire [44:0] buf_acc_data_2_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_5_56_46_sva_mx0;
  wire buf_acc_data_15_11_0_sva_mx0;
  wire [44:0] buf_acc_data_15_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_11_56_46_sva_mx0;
  wire buf_acc_data_2_6_0_sva_mx0;
  wire [44:0] buf_acc_data_2_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_6_56_46_sva_mx0;
  wire buf_acc_data_15_10_0_sva_mx0;
  wire [44:0] buf_acc_data_15_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_10_56_46_sva_mx0;
  wire buf_acc_data_2_7_0_sva_mx0;
  wire [44:0] buf_acc_data_2_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_7_56_46_sva_mx0;
  wire buf_acc_data_15_9_0_sva_mx0;
  wire [44:0] buf_acc_data_15_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_9_56_46_sva_mx0;
  wire buf_acc_data_2_8_0_sva_mx0;
  wire [44:0] buf_acc_data_2_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_8_56_46_sva_mx0;
  wire buf_acc_data_15_8_0_sva_mx0;
  wire [44:0] buf_acc_data_15_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_8_56_46_sva_mx0;
  wire buf_acc_data_2_9_0_sva_mx0;
  wire [44:0] buf_acc_data_2_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_9_56_46_sva_mx0;
  wire buf_acc_data_15_7_0_sva_mx0;
  wire [44:0] buf_acc_data_15_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_7_56_46_sva_mx0;
  wire buf_acc_data_2_10_0_sva_mx0;
  wire [44:0] buf_acc_data_2_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_10_56_46_sva_mx0;
  wire buf_acc_data_15_6_0_sva_mx0;
  wire [44:0] buf_acc_data_15_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_6_56_46_sva_mx0;
  wire buf_acc_data_2_11_0_sva_mx0;
  wire [44:0] buf_acc_data_2_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_11_56_46_sva_mx0;
  wire buf_acc_data_15_5_0_sva_mx0;
  wire [44:0] buf_acc_data_15_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_5_56_46_sva_mx0;
  wire buf_acc_data_2_12_0_sva_mx0;
  wire [44:0] buf_acc_data_2_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_12_56_46_sva_mx0;
  wire buf_acc_data_15_4_0_sva_mx0;
  wire [44:0] buf_acc_data_15_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_4_56_46_sva_mx0;
  wire buf_acc_data_2_13_0_sva_mx0;
  wire [44:0] buf_acc_data_2_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_13_56_46_sva_mx0;
  wire buf_acc_data_15_3_0_sva_mx0;
  wire [44:0] buf_acc_data_15_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_3_56_46_sva_mx0;
  wire buf_acc_data_2_14_0_sva_mx0;
  wire [44:0] buf_acc_data_2_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_14_56_46_sva_mx0;
  wire buf_acc_data_15_2_0_sva_mx0;
  wire [44:0] buf_acc_data_15_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_2_56_46_sva_mx0;
  wire buf_acc_data_2_15_0_sva_mx0;
  wire [44:0] buf_acc_data_2_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_15_56_46_sva_mx0;
  wire buf_acc_data_15_1_0_sva_mx0;
  wire [44:0] buf_acc_data_15_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_1_56_46_sva_mx0;
  wire buf_acc_data_2_16_0_sva_mx0;
  wire [44:0] buf_acc_data_2_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_16_56_46_sva_mx0;
  wire buf_acc_data_15_0_0_sva_mx0;
  wire [44:0] buf_acc_data_15_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_15_0_56_46_sva_mx0;
  wire buf_acc_data_2_17_0_sva_mx0;
  wire [44:0] buf_acc_data_2_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_2_17_56_46_sva_mx0;
  wire buf_acc_data_14_17_0_sva_mx0;
  wire [44:0] buf_acc_data_14_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_17_56_46_sva_mx0;
  wire buf_acc_data_3_0_0_sva_mx0;
  wire [44:0] buf_acc_data_3_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_0_56_46_sva_mx0;
  wire buf_acc_data_14_16_0_sva_mx0;
  wire [44:0] buf_acc_data_14_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_16_56_46_sva_mx0;
  wire buf_acc_data_3_1_0_sva_mx0;
  wire [44:0] buf_acc_data_3_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_1_56_46_sva_mx0;
  wire buf_acc_data_14_15_0_sva_mx0;
  wire [44:0] buf_acc_data_14_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_15_56_46_sva_mx0;
  wire buf_acc_data_3_2_0_sva_mx0;
  wire [44:0] buf_acc_data_3_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_2_56_46_sva_mx0;
  wire buf_acc_data_14_14_0_sva_mx0;
  wire [44:0] buf_acc_data_14_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_14_56_46_sva_mx0;
  wire buf_acc_data_3_3_0_sva_mx0;
  wire [44:0] buf_acc_data_3_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_3_56_46_sva_mx0;
  wire buf_acc_data_14_13_0_sva_mx0;
  wire [44:0] buf_acc_data_14_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_13_56_46_sva_mx0;
  wire buf_acc_data_3_4_0_sva_mx0;
  wire [44:0] buf_acc_data_3_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_4_56_46_sva_mx0;
  wire buf_acc_data_14_12_0_sva_mx0;
  wire [44:0] buf_acc_data_14_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_12_56_46_sva_mx0;
  wire buf_acc_data_3_5_0_sva_mx0;
  wire [44:0] buf_acc_data_3_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_5_56_46_sva_mx0;
  wire buf_acc_data_14_11_0_sva_mx0;
  wire [44:0] buf_acc_data_14_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_11_56_46_sva_mx0;
  wire buf_acc_data_3_6_0_sva_mx0;
  wire [44:0] buf_acc_data_3_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_6_56_46_sva_mx0;
  wire buf_acc_data_14_10_0_sva_mx0;
  wire [44:0] buf_acc_data_14_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_10_56_46_sva_mx0;
  wire buf_acc_data_3_7_0_sva_mx0;
  wire [44:0] buf_acc_data_3_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_7_56_46_sva_mx0;
  wire buf_acc_data_14_9_0_sva_mx0;
  wire [44:0] buf_acc_data_14_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_9_56_46_sva_mx0;
  wire buf_acc_data_3_8_0_sva_mx0;
  wire [44:0] buf_acc_data_3_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_8_56_46_sva_mx0;
  wire buf_acc_data_14_8_0_sva_mx0;
  wire [44:0] buf_acc_data_14_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_8_56_46_sva_mx0;
  wire buf_acc_data_3_9_0_sva_mx0;
  wire [44:0] buf_acc_data_3_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_9_56_46_sva_mx0;
  wire buf_acc_data_14_7_0_sva_mx0;
  wire [44:0] buf_acc_data_14_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_7_56_46_sva_mx0;
  wire buf_acc_data_3_10_0_sva_mx0;
  wire [44:0] buf_acc_data_3_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_10_56_46_sva_mx0;
  wire buf_acc_data_14_6_0_sva_mx0;
  wire [44:0] buf_acc_data_14_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_6_56_46_sva_mx0;
  wire buf_acc_data_3_11_0_sva_mx0;
  wire [44:0] buf_acc_data_3_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_11_56_46_sva_mx0;
  wire buf_acc_data_14_5_0_sva_mx0;
  wire [44:0] buf_acc_data_14_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_5_56_46_sva_mx0;
  wire buf_acc_data_3_12_0_sva_mx0;
  wire [44:0] buf_acc_data_3_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_12_56_46_sva_mx0;
  wire buf_acc_data_14_4_0_sva_mx0;
  wire [44:0] buf_acc_data_14_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_4_56_46_sva_mx0;
  wire buf_acc_data_3_13_0_sva_mx0;
  wire [44:0] buf_acc_data_3_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_13_56_46_sva_mx0;
  wire buf_acc_data_14_3_0_sva_mx0;
  wire [44:0] buf_acc_data_14_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_3_56_46_sva_mx0;
  wire buf_acc_data_3_14_0_sva_mx0;
  wire [44:0] buf_acc_data_3_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_14_56_46_sva_mx0;
  wire buf_acc_data_14_2_0_sva_mx0;
  wire [44:0] buf_acc_data_14_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_2_56_46_sva_mx0;
  wire buf_acc_data_3_15_0_sva_mx0;
  wire [44:0] buf_acc_data_3_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_15_56_46_sva_mx0;
  wire buf_acc_data_14_1_0_sva_mx0;
  wire [44:0] buf_acc_data_14_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_1_56_46_sva_mx0;
  wire buf_acc_data_3_16_0_sva_mx0;
  wire [44:0] buf_acc_data_3_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_16_56_46_sva_mx0;
  wire buf_acc_data_14_0_0_sva_mx0;
  wire [44:0] buf_acc_data_14_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_14_0_56_46_sva_mx0;
  wire buf_acc_data_3_17_0_sva_mx0;
  wire [44:0] buf_acc_data_3_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_3_17_56_46_sva_mx0;
  wire buf_acc_data_13_17_0_sva_mx0;
  wire [44:0] buf_acc_data_13_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_17_56_46_sva_mx0;
  wire buf_acc_data_4_0_0_sva_mx0;
  wire [44:0] buf_acc_data_4_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_0_56_46_sva_mx0;
  wire buf_acc_data_13_16_0_sva_mx0;
  wire [44:0] buf_acc_data_13_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_16_56_46_sva_mx0;
  wire buf_acc_data_4_1_0_sva_mx0;
  wire [44:0] buf_acc_data_4_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_1_56_46_sva_mx0;
  wire buf_acc_data_13_15_0_sva_mx0;
  wire [44:0] buf_acc_data_13_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_15_56_46_sva_mx0;
  wire buf_acc_data_4_2_0_sva_mx0;
  wire [44:0] buf_acc_data_4_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_2_56_46_sva_mx0;
  wire buf_acc_data_13_14_0_sva_mx0;
  wire [44:0] buf_acc_data_13_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_14_56_46_sva_mx0;
  wire buf_acc_data_4_3_0_sva_mx0;
  wire [44:0] buf_acc_data_4_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_3_56_46_sva_mx0;
  wire buf_acc_data_13_13_0_sva_mx0;
  wire [44:0] buf_acc_data_13_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_13_56_46_sva_mx0;
  wire buf_acc_data_4_4_0_sva_mx0;
  wire [44:0] buf_acc_data_4_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_4_56_46_sva_mx0;
  wire buf_acc_data_13_12_0_sva_mx0;
  wire [44:0] buf_acc_data_13_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_12_56_46_sva_mx0;
  wire buf_acc_data_4_5_0_sva_mx0;
  wire [44:0] buf_acc_data_4_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_5_56_46_sva_mx0;
  wire buf_acc_data_13_11_0_sva_mx0;
  wire [44:0] buf_acc_data_13_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_11_56_46_sva_mx0;
  wire buf_acc_data_4_6_0_sva_mx0;
  wire [44:0] buf_acc_data_4_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_6_56_46_sva_mx0;
  wire buf_acc_data_13_10_0_sva_mx0;
  wire [44:0] buf_acc_data_13_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_10_56_46_sva_mx0;
  wire buf_acc_data_4_7_0_sva_mx0;
  wire [44:0] buf_acc_data_4_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_7_56_46_sva_mx0;
  wire buf_acc_data_13_9_0_sva_mx0;
  wire [44:0] buf_acc_data_13_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_9_56_46_sva_mx0;
  wire buf_acc_data_4_8_0_sva_mx0;
  wire [44:0] buf_acc_data_4_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_8_56_46_sva_mx0;
  wire buf_acc_data_13_8_0_sva_mx0;
  wire [44:0] buf_acc_data_13_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_8_56_46_sva_mx0;
  wire buf_acc_data_4_9_0_sva_mx0;
  wire [44:0] buf_acc_data_4_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_9_56_46_sva_mx0;
  wire buf_acc_data_13_7_0_sva_mx0;
  wire [44:0] buf_acc_data_13_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_7_56_46_sva_mx0;
  wire buf_acc_data_4_10_0_sva_mx0;
  wire [44:0] buf_acc_data_4_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_10_56_46_sva_mx0;
  wire buf_acc_data_13_6_0_sva_mx0;
  wire [44:0] buf_acc_data_13_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_6_56_46_sva_mx0;
  wire buf_acc_data_4_11_0_sva_mx0;
  wire [44:0] buf_acc_data_4_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_11_56_46_sva_mx0;
  wire buf_acc_data_13_5_0_sva_mx0;
  wire [44:0] buf_acc_data_13_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_5_56_46_sva_mx0;
  wire buf_acc_data_4_12_0_sva_mx0;
  wire [44:0] buf_acc_data_4_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_12_56_46_sva_mx0;
  wire buf_acc_data_13_4_0_sva_mx0;
  wire [44:0] buf_acc_data_13_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_4_56_46_sva_mx0;
  wire buf_acc_data_4_13_0_sva_mx0;
  wire [44:0] buf_acc_data_4_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_13_56_46_sva_mx0;
  wire buf_acc_data_13_3_0_sva_mx0;
  wire [44:0] buf_acc_data_13_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_3_56_46_sva_mx0;
  wire buf_acc_data_4_14_0_sva_mx0;
  wire [44:0] buf_acc_data_4_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_14_56_46_sva_mx0;
  wire buf_acc_data_13_2_0_sva_mx0;
  wire [44:0] buf_acc_data_13_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_2_56_46_sva_mx0;
  wire buf_acc_data_4_15_0_sva_mx0;
  wire [44:0] buf_acc_data_4_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_15_56_46_sva_mx0;
  wire buf_acc_data_13_1_0_sva_mx0;
  wire [44:0] buf_acc_data_13_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_1_56_46_sva_mx0;
  wire buf_acc_data_4_16_0_sva_mx0;
  wire [44:0] buf_acc_data_4_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_16_56_46_sva_mx0;
  wire buf_acc_data_13_0_0_sva_mx0;
  wire [44:0] buf_acc_data_13_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_13_0_56_46_sva_mx0;
  wire buf_acc_data_4_17_0_sva_mx0;
  wire [44:0] buf_acc_data_4_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_4_17_56_46_sva_mx0;
  wire buf_acc_data_12_17_0_sva_mx0;
  wire [44:0] buf_acc_data_12_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_17_56_46_sva_mx0;
  wire buf_acc_data_5_0_0_sva_mx0;
  wire [44:0] buf_acc_data_5_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_0_56_46_sva_mx0;
  wire buf_acc_data_12_16_0_sva_mx0;
  wire [44:0] buf_acc_data_12_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_16_56_46_sva_mx0;
  wire buf_acc_data_5_1_0_sva_mx0;
  wire [44:0] buf_acc_data_5_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_1_56_46_sva_mx0;
  wire buf_acc_data_12_15_0_sva_mx0;
  wire [44:0] buf_acc_data_12_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_15_56_46_sva_mx0;
  wire buf_acc_data_5_2_0_sva_mx0;
  wire [44:0] buf_acc_data_5_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_2_56_46_sva_mx0;
  wire buf_acc_data_12_14_0_sva_mx0;
  wire [44:0] buf_acc_data_12_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_14_56_46_sva_mx0;
  wire buf_acc_data_5_3_0_sva_mx0;
  wire [44:0] buf_acc_data_5_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_3_56_46_sva_mx0;
  wire buf_acc_data_12_13_0_sva_mx0;
  wire [44:0] buf_acc_data_12_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_13_56_46_sva_mx0;
  wire buf_acc_data_5_4_0_sva_mx0;
  wire [44:0] buf_acc_data_5_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_4_56_46_sva_mx0;
  wire buf_acc_data_12_12_0_sva_mx0;
  wire [44:0] buf_acc_data_12_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_12_56_46_sva_mx0;
  wire buf_acc_data_5_5_0_sva_mx0;
  wire [44:0] buf_acc_data_5_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_5_56_46_sva_mx0;
  wire buf_acc_data_12_11_0_sva_mx0;
  wire [44:0] buf_acc_data_12_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_11_56_46_sva_mx0;
  wire buf_acc_data_5_6_0_sva_mx0;
  wire [44:0] buf_acc_data_5_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_6_56_46_sva_mx0;
  wire buf_acc_data_12_10_0_sva_mx0;
  wire [44:0] buf_acc_data_12_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_10_56_46_sva_mx0;
  wire buf_acc_data_5_7_0_sva_mx0;
  wire [44:0] buf_acc_data_5_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_7_56_46_sva_mx0;
  wire buf_acc_data_12_9_0_sva_mx0;
  wire [44:0] buf_acc_data_12_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_9_56_46_sva_mx0;
  wire buf_acc_data_5_8_0_sva_mx0;
  wire [44:0] buf_acc_data_5_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_8_56_46_sva_mx0;
  wire buf_acc_data_12_8_0_sva_mx0;
  wire [44:0] buf_acc_data_12_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_8_56_46_sva_mx0;
  wire buf_acc_data_5_9_0_sva_mx0;
  wire [44:0] buf_acc_data_5_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_9_56_46_sva_mx0;
  wire buf_acc_data_12_7_0_sva_mx0;
  wire [44:0] buf_acc_data_12_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_7_56_46_sva_mx0;
  wire buf_acc_data_5_10_0_sva_mx0;
  wire [44:0] buf_acc_data_5_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_10_56_46_sva_mx0;
  wire buf_acc_data_12_6_0_sva_mx0;
  wire [44:0] buf_acc_data_12_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_6_56_46_sva_mx0;
  wire buf_acc_data_5_11_0_sva_mx0;
  wire [44:0] buf_acc_data_5_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_11_56_46_sva_mx0;
  wire buf_acc_data_12_5_0_sva_mx0;
  wire [44:0] buf_acc_data_12_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_5_56_46_sva_mx0;
  wire buf_acc_data_5_12_0_sva_mx0;
  wire [44:0] buf_acc_data_5_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_12_56_46_sva_mx0;
  wire buf_acc_data_12_4_0_sva_mx0;
  wire [44:0] buf_acc_data_12_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_4_56_46_sva_mx0;
  wire buf_acc_data_5_13_0_sva_mx0;
  wire [44:0] buf_acc_data_5_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_13_56_46_sva_mx0;
  wire buf_acc_data_12_3_0_sva_mx0;
  wire [44:0] buf_acc_data_12_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_3_56_46_sva_mx0;
  wire buf_acc_data_5_14_0_sva_mx0;
  wire [44:0] buf_acc_data_5_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_14_56_46_sva_mx0;
  wire buf_acc_data_12_2_0_sva_mx0;
  wire [44:0] buf_acc_data_12_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_2_56_46_sva_mx0;
  wire buf_acc_data_5_15_0_sva_mx0;
  wire [44:0] buf_acc_data_5_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_15_56_46_sva_mx0;
  wire buf_acc_data_12_1_0_sva_mx0;
  wire [44:0] buf_acc_data_12_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_1_56_46_sva_mx0;
  wire buf_acc_data_5_16_0_sva_mx0;
  wire [44:0] buf_acc_data_5_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_16_56_46_sva_mx0;
  wire buf_acc_data_12_0_0_sva_mx0;
  wire [44:0] buf_acc_data_12_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_12_0_56_46_sva_mx0;
  wire buf_acc_data_5_17_0_sva_mx0;
  wire [44:0] buf_acc_data_5_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_5_17_56_46_sva_mx0;
  wire buf_acc_data_11_17_0_sva_mx0;
  wire [44:0] buf_acc_data_11_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_17_56_46_sva_mx0;
  wire buf_acc_data_6_0_0_sva_mx0;
  wire [44:0] buf_acc_data_6_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_0_56_46_sva_mx0;
  wire buf_acc_data_11_16_0_sva_mx0;
  wire [44:0] buf_acc_data_11_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_16_56_46_sva_mx0;
  wire buf_acc_data_6_1_0_sva_mx0;
  wire [44:0] buf_acc_data_6_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_1_56_46_sva_mx0;
  wire buf_acc_data_11_15_0_sva_mx0;
  wire [44:0] buf_acc_data_11_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_15_56_46_sva_mx0;
  wire buf_acc_data_6_2_0_sva_mx0;
  wire [44:0] buf_acc_data_6_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_2_56_46_sva_mx0;
  wire buf_acc_data_11_14_0_sva_mx0;
  wire [44:0] buf_acc_data_11_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_14_56_46_sva_mx0;
  wire buf_acc_data_6_3_0_sva_mx0;
  wire [44:0] buf_acc_data_6_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_3_56_46_sva_mx0;
  wire buf_acc_data_11_13_0_sva_mx0;
  wire [44:0] buf_acc_data_11_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_13_56_46_sva_mx0;
  wire buf_acc_data_6_4_0_sva_mx0;
  wire [44:0] buf_acc_data_6_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_4_56_46_sva_mx0;
  wire buf_acc_data_11_12_0_sva_mx0;
  wire [44:0] buf_acc_data_11_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_12_56_46_sva_mx0;
  wire buf_acc_data_6_5_0_sva_mx0;
  wire [44:0] buf_acc_data_6_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_5_56_46_sva_mx0;
  wire buf_acc_data_11_11_0_sva_mx0;
  wire [44:0] buf_acc_data_11_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_11_56_46_sva_mx0;
  wire buf_acc_data_6_6_0_sva_mx0;
  wire [44:0] buf_acc_data_6_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_6_56_46_sva_mx0;
  wire buf_acc_data_11_10_0_sva_mx0;
  wire [44:0] buf_acc_data_11_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_10_56_46_sva_mx0;
  wire buf_acc_data_6_7_0_sva_mx0;
  wire [44:0] buf_acc_data_6_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_7_56_46_sva_mx0;
  wire buf_acc_data_11_9_0_sva_mx0;
  wire [44:0] buf_acc_data_11_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_9_56_46_sva_mx0;
  wire buf_acc_data_6_8_0_sva_mx0;
  wire [44:0] buf_acc_data_6_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_8_56_46_sva_mx0;
  wire buf_acc_data_11_8_0_sva_mx0;
  wire [44:0] buf_acc_data_11_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_8_56_46_sva_mx0;
  wire buf_acc_data_6_9_0_sva_mx0;
  wire [44:0] buf_acc_data_6_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_9_56_46_sva_mx0;
  wire buf_acc_data_11_7_0_sva_mx0;
  wire [44:0] buf_acc_data_11_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_7_56_46_sva_mx0;
  wire buf_acc_data_6_10_0_sva_mx0;
  wire [44:0] buf_acc_data_6_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_10_56_46_sva_mx0;
  wire buf_acc_data_11_6_0_sva_mx0;
  wire [44:0] buf_acc_data_11_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_6_56_46_sva_mx0;
  wire buf_acc_data_6_11_0_sva_mx0;
  wire [44:0] buf_acc_data_6_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_11_56_46_sva_mx0;
  wire buf_acc_data_11_5_0_sva_mx0;
  wire [44:0] buf_acc_data_11_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_5_56_46_sva_mx0;
  wire buf_acc_data_6_12_0_sva_mx0;
  wire [44:0] buf_acc_data_6_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_12_56_46_sva_mx0;
  wire buf_acc_data_11_4_0_sva_mx0;
  wire [44:0] buf_acc_data_11_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_4_56_46_sva_mx0;
  wire buf_acc_data_6_13_0_sva_mx0;
  wire [44:0] buf_acc_data_6_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_13_56_46_sva_mx0;
  wire buf_acc_data_11_3_0_sva_mx0;
  wire [44:0] buf_acc_data_11_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_3_56_46_sva_mx0;
  wire buf_acc_data_6_14_0_sva_mx0;
  wire [44:0] buf_acc_data_6_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_14_56_46_sva_mx0;
  wire buf_acc_data_11_2_0_sva_mx0;
  wire [44:0] buf_acc_data_11_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_2_56_46_sva_mx0;
  wire buf_acc_data_6_15_0_sva_mx0;
  wire [44:0] buf_acc_data_6_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_15_56_46_sva_mx0;
  wire buf_acc_data_11_1_0_sva_mx0;
  wire [44:0] buf_acc_data_11_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_1_56_46_sva_mx0;
  wire buf_acc_data_6_16_0_sva_mx0;
  wire [44:0] buf_acc_data_6_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_16_56_46_sva_mx0;
  wire buf_acc_data_11_0_0_sva_mx0;
  wire [44:0] buf_acc_data_11_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_11_0_56_46_sva_mx0;
  wire buf_acc_data_6_17_0_sva_mx0;
  wire [44:0] buf_acc_data_6_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_6_17_56_46_sva_mx0;
  wire buf_acc_data_10_17_0_sva_mx0;
  wire [44:0] buf_acc_data_10_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_17_56_46_sva_mx0;
  wire buf_acc_data_7_0_0_sva_mx0;
  wire [44:0] buf_acc_data_7_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_0_56_46_sva_mx0;
  wire buf_acc_data_10_16_0_sva_mx0;
  wire [44:0] buf_acc_data_10_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_16_56_46_sva_mx0;
  wire buf_acc_data_7_1_0_sva_mx0;
  wire [44:0] buf_acc_data_7_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_1_56_46_sva_mx0;
  wire buf_acc_data_10_15_0_sva_mx0;
  wire [44:0] buf_acc_data_10_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_15_56_46_sva_mx0;
  wire buf_acc_data_7_2_0_sva_mx0;
  wire [44:0] buf_acc_data_7_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_2_56_46_sva_mx0;
  wire buf_acc_data_10_14_0_sva_mx0;
  wire [44:0] buf_acc_data_10_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_14_56_46_sva_mx0;
  wire buf_acc_data_7_3_0_sva_mx0;
  wire [44:0] buf_acc_data_7_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_3_56_46_sva_mx0;
  wire buf_acc_data_10_13_0_sva_mx0;
  wire [44:0] buf_acc_data_10_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_13_56_46_sva_mx0;
  wire buf_acc_data_7_4_0_sva_mx0;
  wire [44:0] buf_acc_data_7_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_4_56_46_sva_mx0;
  wire buf_acc_data_10_12_0_sva_mx0;
  wire [44:0] buf_acc_data_10_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_12_56_46_sva_mx0;
  wire buf_acc_data_7_5_0_sva_mx0;
  wire [44:0] buf_acc_data_7_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_5_56_46_sva_mx0;
  wire buf_acc_data_10_11_0_sva_mx0;
  wire [44:0] buf_acc_data_10_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_11_56_46_sva_mx0;
  wire buf_acc_data_7_6_0_sva_mx0;
  wire [44:0] buf_acc_data_7_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_6_56_46_sva_mx0;
  wire buf_acc_data_10_10_0_sva_mx0;
  wire [44:0] buf_acc_data_10_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_10_56_46_sva_mx0;
  wire buf_acc_data_7_7_0_sva_mx0;
  wire [44:0] buf_acc_data_7_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_7_56_46_sva_mx0;
  wire buf_acc_data_10_9_0_sva_mx0;
  wire [44:0] buf_acc_data_10_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_9_56_46_sva_mx0;
  wire buf_acc_data_7_8_0_sva_mx0;
  wire [44:0] buf_acc_data_7_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_8_56_46_sva_mx0;
  wire buf_acc_data_10_8_0_sva_mx0;
  wire [44:0] buf_acc_data_10_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_8_56_46_sva_mx0;
  wire buf_acc_data_7_9_0_sva_mx0;
  wire [44:0] buf_acc_data_7_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_9_56_46_sva_mx0;
  wire buf_acc_data_10_7_0_sva_mx0;
  wire [44:0] buf_acc_data_10_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_7_56_46_sva_mx0;
  wire buf_acc_data_7_10_0_sva_mx0;
  wire [44:0] buf_acc_data_7_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_10_56_46_sva_mx0;
  wire buf_acc_data_10_6_0_sva_mx0;
  wire [44:0] buf_acc_data_10_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_6_56_46_sva_mx0;
  wire buf_acc_data_7_11_0_sva_mx0;
  wire [44:0] buf_acc_data_7_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_11_56_46_sva_mx0;
  wire buf_acc_data_10_5_0_sva_mx0;
  wire [44:0] buf_acc_data_10_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_5_56_46_sva_mx0;
  wire buf_acc_data_7_12_0_sva_mx0;
  wire [44:0] buf_acc_data_7_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_12_56_46_sva_mx0;
  wire buf_acc_data_10_4_0_sva_mx0;
  wire [44:0] buf_acc_data_10_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_4_56_46_sva_mx0;
  wire buf_acc_data_7_13_0_sva_mx0;
  wire [44:0] buf_acc_data_7_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_13_56_46_sva_mx0;
  wire buf_acc_data_10_3_0_sva_mx0;
  wire [44:0] buf_acc_data_10_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_3_56_46_sva_mx0;
  wire buf_acc_data_7_14_0_sva_mx0;
  wire [44:0] buf_acc_data_7_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_14_56_46_sva_mx0;
  wire buf_acc_data_10_2_0_sva_mx0;
  wire [44:0] buf_acc_data_10_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_2_56_46_sva_mx0;
  wire buf_acc_data_7_15_0_sva_mx0;
  wire [44:0] buf_acc_data_7_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_15_56_46_sva_mx0;
  wire buf_acc_data_10_1_0_sva_mx0;
  wire [44:0] buf_acc_data_10_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_1_56_46_sva_mx0;
  wire buf_acc_data_7_16_0_sva_mx0;
  wire [44:0] buf_acc_data_7_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_16_56_46_sva_mx0;
  wire buf_acc_data_10_0_0_sva_mx0;
  wire [44:0] buf_acc_data_10_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_10_0_56_46_sva_mx0;
  wire buf_acc_data_7_17_0_sva_mx0;
  wire [44:0] buf_acc_data_7_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_7_17_56_46_sva_mx0;
  wire buf_acc_data_9_17_0_sva_mx0;
  wire [44:0] buf_acc_data_9_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_17_56_46_sva_mx0;
  wire buf_acc_data_8_0_0_sva_mx0;
  wire [44:0] buf_acc_data_8_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_0_56_46_sva_mx0;
  wire buf_acc_data_9_16_0_sva_mx0;
  wire [44:0] buf_acc_data_9_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_16_56_46_sva_mx0;
  wire buf_acc_data_8_1_0_sva_mx0;
  wire [44:0] buf_acc_data_8_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_1_56_46_sva_mx0;
  wire buf_acc_data_9_15_0_sva_mx0;
  wire [44:0] buf_acc_data_9_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_15_56_46_sva_mx0;
  wire buf_acc_data_8_2_0_sva_mx0;
  wire [44:0] buf_acc_data_8_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_2_56_46_sva_mx0;
  wire buf_acc_data_9_14_0_sva_mx0;
  wire [44:0] buf_acc_data_9_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_14_56_46_sva_mx0;
  wire buf_acc_data_8_3_0_sva_mx0;
  wire [44:0] buf_acc_data_8_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_3_56_46_sva_mx0;
  wire buf_acc_data_9_13_0_sva_mx0;
  wire [44:0] buf_acc_data_9_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_13_56_46_sva_mx0;
  wire buf_acc_data_8_4_0_sva_mx0;
  wire [44:0] buf_acc_data_8_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_4_56_46_sva_mx0;
  wire buf_acc_data_9_12_0_sva_mx0;
  wire [44:0] buf_acc_data_9_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_12_56_46_sva_mx0;
  wire buf_acc_data_8_5_0_sva_mx0;
  wire [44:0] buf_acc_data_8_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_5_56_46_sva_mx0;
  wire buf_acc_data_9_11_0_sva_mx0;
  wire [44:0] buf_acc_data_9_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_11_56_46_sva_mx0;
  wire buf_acc_data_8_6_0_sva_mx0;
  wire [44:0] buf_acc_data_8_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_6_56_46_sva_mx0;
  wire buf_acc_data_9_10_0_sva_mx0;
  wire [44:0] buf_acc_data_9_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_10_56_46_sva_mx0;
  wire buf_acc_data_8_7_0_sva_mx0;
  wire [44:0] buf_acc_data_8_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_7_56_46_sva_mx0;
  wire buf_acc_data_9_9_0_sva_mx0;
  wire [44:0] buf_acc_data_9_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_9_56_46_sva_mx0;
  wire buf_acc_data_8_8_0_sva_mx0;
  wire [44:0] buf_acc_data_8_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_8_56_46_sva_mx0;
  wire buf_acc_data_9_8_0_sva_mx0;
  wire [44:0] buf_acc_data_9_8_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_8_56_46_sva_mx0;
  wire buf_acc_data_8_9_0_sva_mx0;
  wire [44:0] buf_acc_data_8_9_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_9_56_46_sva_mx0;
  wire buf_acc_data_9_7_0_sva_mx0;
  wire [44:0] buf_acc_data_9_7_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_7_56_46_sva_mx0;
  wire buf_acc_data_8_10_0_sva_mx0;
  wire [44:0] buf_acc_data_8_10_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_10_56_46_sva_mx0;
  wire buf_acc_data_9_6_0_sva_mx0;
  wire [44:0] buf_acc_data_9_6_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_6_56_46_sva_mx0;
  wire buf_acc_data_8_11_0_sva_mx0;
  wire [44:0] buf_acc_data_8_11_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_11_56_46_sva_mx0;
  wire buf_acc_data_9_5_0_sva_mx0;
  wire [44:0] buf_acc_data_9_5_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_5_56_46_sva_mx0;
  wire buf_acc_data_8_12_0_sva_mx0;
  wire [44:0] buf_acc_data_8_12_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_12_56_46_sva_mx0;
  wire buf_acc_data_9_4_0_sva_mx0;
  wire [44:0] buf_acc_data_9_4_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_4_56_46_sva_mx0;
  wire buf_acc_data_8_13_0_sva_mx0;
  wire [44:0] buf_acc_data_8_13_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_13_56_46_sva_mx0;
  wire buf_acc_data_9_3_0_sva_mx0;
  wire [44:0] buf_acc_data_9_3_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_3_56_46_sva_mx0;
  wire buf_acc_data_8_14_0_sva_mx0;
  wire [44:0] buf_acc_data_8_14_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_14_56_46_sva_mx0;
  wire buf_acc_data_9_2_0_sva_mx0;
  wire [44:0] buf_acc_data_9_2_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_2_56_46_sva_mx0;
  wire buf_acc_data_8_15_0_sva_mx0;
  wire [44:0] buf_acc_data_8_15_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_15_56_46_sva_mx0;
  wire buf_acc_data_9_1_0_sva_mx0;
  wire [44:0] buf_acc_data_9_1_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_1_56_46_sva_mx0;
  wire buf_acc_data_8_16_0_sva_mx0;
  wire [44:0] buf_acc_data_8_16_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_16_56_46_sva_mx0;
  wire buf_acc_data_9_0_0_sva_mx0;
  wire [44:0] buf_acc_data_9_0_45_1_sva_mx0;
  wire [10:0] buf_acc_data_9_0_56_46_sva_mx0;
  wire buf_acc_data_8_17_0_sva_mx0;
  wire [44:0] buf_acc_data_8_17_45_1_sva_mx0;
  wire [10:0] buf_acc_data_8_17_56_46_sva_mx0;
  wire CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_mx1;
  wire CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_mx1;
  wire CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1;
  wire buf_acc_data_0_0_0_sva_dfm_mx0;
  wire buf_acc_data_0_1_0_sva_dfm_mx0;
  wire buf_acc_data_0_2_0_sva_dfm_mx0;
  wire buf_acc_data_0_3_0_sva_dfm_mx0;
  wire buf_acc_data_0_4_0_sva_dfm_mx0;
  wire buf_acc_data_0_5_0_sva_dfm_mx0;
  wire buf_acc_data_0_6_0_sva_dfm_mx0;
  wire buf_acc_data_0_7_0_sva_dfm_mx0;
  wire buf_acc_data_0_8_0_sva_dfm_mx0;
  wire buf_acc_data_0_9_0_sva_dfm_mx0;
  wire buf_acc_data_0_10_0_sva_dfm_mx0;
  wire buf_acc_data_0_11_0_sva_dfm_mx0;
  wire buf_acc_data_0_12_0_sva_dfm_mx0;
  wire buf_acc_data_0_13_0_sva_dfm_mx0;
  wire buf_acc_data_0_14_0_sva_dfm_mx0;
  wire buf_acc_data_0_15_0_sva_dfm_mx0;
  wire buf_acc_data_0_16_0_sva_dfm_mx0;
  wire buf_acc_data_0_17_0_sva_dfm_mx0;
  wire buf_acc_data_1_0_0_sva_dfm_mx0;
  wire buf_acc_data_1_1_0_sva_dfm_mx0;
  wire buf_acc_data_1_2_0_sva_dfm_mx0;
  wire buf_acc_data_1_3_0_sva_dfm_mx0;
  wire buf_acc_data_1_4_0_sva_dfm_mx0;
  wire buf_acc_data_1_5_0_sva_dfm_mx0;
  wire buf_acc_data_1_6_0_sva_dfm_mx0;
  wire buf_acc_data_1_7_0_sva_dfm_mx0;
  wire buf_acc_data_1_8_0_sva_dfm_mx0;
  wire buf_acc_data_1_9_0_sva_dfm_mx0;
  wire buf_acc_data_1_10_0_sva_dfm_mx0;
  wire buf_acc_data_1_11_0_sva_dfm_mx0;
  wire buf_acc_data_1_12_0_sva_dfm_mx0;
  wire buf_acc_data_1_13_0_sva_dfm_mx0;
  wire buf_acc_data_1_14_0_sva_dfm_mx0;
  wire buf_acc_data_1_15_0_sva_dfm_mx0;
  wire buf_acc_data_1_16_0_sva_dfm_mx0;
  wire buf_acc_data_1_17_0_sva_dfm_mx0;
  wire buf_acc_data_2_0_0_sva_dfm_mx0;
  wire buf_acc_data_2_1_0_sva_dfm_mx0;
  wire buf_acc_data_2_2_0_sva_dfm_mx0;
  wire buf_acc_data_2_3_0_sva_dfm_mx0;
  wire buf_acc_data_2_4_0_sva_dfm_mx0;
  wire buf_acc_data_2_5_0_sva_dfm_mx0;
  wire buf_acc_data_2_6_0_sva_dfm_mx0;
  wire buf_acc_data_2_7_0_sva_dfm_mx0;
  wire buf_acc_data_2_8_0_sva_dfm_mx0;
  wire buf_acc_data_2_9_0_sva_dfm_mx0;
  wire buf_acc_data_2_10_0_sva_dfm_mx0;
  wire buf_acc_data_2_11_0_sva_dfm_mx0;
  wire buf_acc_data_2_12_0_sva_dfm_mx0;
  wire buf_acc_data_2_13_0_sva_dfm_mx0;
  wire buf_acc_data_2_14_0_sva_dfm_mx0;
  wire buf_acc_data_2_15_0_sva_dfm_mx0;
  wire buf_acc_data_2_16_0_sva_dfm_mx0;
  wire buf_acc_data_2_17_0_sva_dfm_mx0;
  wire buf_acc_data_3_0_0_sva_dfm_mx0;
  wire buf_acc_data_3_1_0_sva_dfm_mx0;
  wire buf_acc_data_3_2_0_sva_dfm_mx0;
  wire buf_acc_data_3_3_0_sva_dfm_mx0;
  wire buf_acc_data_3_4_0_sva_dfm_mx0;
  wire buf_acc_data_3_5_0_sva_dfm_mx0;
  wire buf_acc_data_3_6_0_sva_dfm_mx0;
  wire buf_acc_data_3_7_0_sva_dfm_mx0;
  wire buf_acc_data_3_8_0_sva_dfm_mx0;
  wire buf_acc_data_3_9_0_sva_dfm_mx0;
  wire buf_acc_data_3_10_0_sva_dfm_mx0;
  wire buf_acc_data_3_11_0_sva_dfm_mx0;
  wire buf_acc_data_3_12_0_sva_dfm_mx0;
  wire buf_acc_data_3_13_0_sva_dfm_mx0;
  wire buf_acc_data_3_14_0_sva_dfm_mx0;
  wire buf_acc_data_3_15_0_sva_dfm_mx0;
  wire buf_acc_data_3_16_0_sva_dfm_mx0;
  wire buf_acc_data_3_17_0_sva_dfm_mx0;
  wire buf_acc_data_4_0_0_sva_dfm_mx0;
  wire buf_acc_data_4_1_0_sva_dfm_mx0;
  wire buf_acc_data_4_2_0_sva_dfm_mx0;
  wire buf_acc_data_4_3_0_sva_dfm_mx0;
  wire buf_acc_data_4_4_0_sva_dfm_mx0;
  wire buf_acc_data_4_5_0_sva_dfm_mx0;
  wire buf_acc_data_4_6_0_sva_dfm_mx0;
  wire buf_acc_data_4_7_0_sva_dfm_mx0;
  wire buf_acc_data_4_8_0_sva_dfm_mx0;
  wire buf_acc_data_4_9_0_sva_dfm_mx0;
  wire buf_acc_data_4_10_0_sva_dfm_mx0;
  wire buf_acc_data_4_11_0_sva_dfm_mx0;
  wire buf_acc_data_4_12_0_sva_dfm_mx0;
  wire buf_acc_data_4_13_0_sva_dfm_mx0;
  wire buf_acc_data_4_14_0_sva_dfm_mx0;
  wire buf_acc_data_4_15_0_sva_dfm_mx0;
  wire buf_acc_data_4_16_0_sva_dfm_mx0;
  wire buf_acc_data_4_17_0_sva_dfm_mx0;
  wire buf_acc_data_5_0_0_sva_dfm_mx0;
  wire buf_acc_data_5_1_0_sva_dfm_mx0;
  wire buf_acc_data_5_2_0_sva_dfm_mx0;
  wire buf_acc_data_5_3_0_sva_dfm_mx0;
  wire buf_acc_data_5_4_0_sva_dfm_mx0;
  wire buf_acc_data_5_5_0_sva_dfm_mx0;
  wire buf_acc_data_5_6_0_sva_dfm_mx0;
  wire buf_acc_data_5_7_0_sva_dfm_mx0;
  wire buf_acc_data_5_8_0_sva_dfm_mx0;
  wire buf_acc_data_5_9_0_sva_dfm_mx0;
  wire buf_acc_data_5_10_0_sva_dfm_mx0;
  wire buf_acc_data_5_11_0_sva_dfm_mx0;
  wire buf_acc_data_5_12_0_sva_dfm_mx0;
  wire buf_acc_data_5_13_0_sva_dfm_mx0;
  wire buf_acc_data_5_14_0_sva_dfm_mx0;
  wire buf_acc_data_5_15_0_sva_dfm_mx0;
  wire buf_acc_data_5_16_0_sva_dfm_mx0;
  wire buf_acc_data_5_17_0_sva_dfm_mx0;
  wire buf_acc_data_6_0_0_sva_dfm_mx0;
  wire buf_acc_data_6_1_0_sva_dfm_mx0;
  wire buf_acc_data_6_2_0_sva_dfm_mx0;
  wire buf_acc_data_6_3_0_sva_dfm_mx0;
  wire buf_acc_data_6_4_0_sva_dfm_mx0;
  wire buf_acc_data_6_5_0_sva_dfm_mx0;
  wire buf_acc_data_6_6_0_sva_dfm_mx0;
  wire buf_acc_data_6_7_0_sva_dfm_mx0;
  wire buf_acc_data_6_8_0_sva_dfm_mx0;
  wire buf_acc_data_6_9_0_sva_dfm_mx0;
  wire buf_acc_data_6_10_0_sva_dfm_mx0;
  wire buf_acc_data_6_11_0_sva_dfm_mx0;
  wire buf_acc_data_6_12_0_sva_dfm_mx0;
  wire buf_acc_data_6_13_0_sva_dfm_mx0;
  wire buf_acc_data_6_14_0_sva_dfm_mx0;
  wire buf_acc_data_6_15_0_sva_dfm_mx0;
  wire buf_acc_data_6_16_0_sva_dfm_mx0;
  wire buf_acc_data_6_17_0_sva_dfm_mx0;
  wire buf_acc_data_7_0_0_sva_dfm_mx0;
  wire buf_acc_data_7_1_0_sva_dfm_mx0;
  wire buf_acc_data_7_2_0_sva_dfm_mx0;
  wire buf_acc_data_7_3_0_sva_dfm_mx0;
  wire buf_acc_data_7_4_0_sva_dfm_mx0;
  wire buf_acc_data_7_5_0_sva_dfm_mx0;
  wire buf_acc_data_7_6_0_sva_dfm_mx0;
  wire buf_acc_data_7_7_0_sva_dfm_mx0;
  wire buf_acc_data_7_8_0_sva_dfm_mx0;
  wire buf_acc_data_7_9_0_sva_dfm_mx0;
  wire buf_acc_data_7_10_0_sva_dfm_mx0;
  wire buf_acc_data_7_11_0_sva_dfm_mx0;
  wire buf_acc_data_7_12_0_sva_dfm_mx0;
  wire buf_acc_data_7_13_0_sva_dfm_mx0;
  wire buf_acc_data_7_14_0_sva_dfm_mx0;
  wire buf_acc_data_7_15_0_sva_dfm_mx0;
  wire buf_acc_data_7_16_0_sva_dfm_mx0;
  wire buf_acc_data_7_17_0_sva_dfm_mx0;
  wire buf_acc_data_8_0_0_sva_dfm_mx0;
  wire buf_acc_data_8_1_0_sva_dfm_mx0;
  wire buf_acc_data_8_2_0_sva_dfm_mx0;
  wire buf_acc_data_8_3_0_sva_dfm_mx0;
  wire buf_acc_data_8_4_0_sva_dfm_mx0;
  wire buf_acc_data_8_5_0_sva_dfm_mx0;
  wire buf_acc_data_8_6_0_sva_dfm_mx0;
  wire buf_acc_data_8_7_0_sva_dfm_mx0;
  wire buf_acc_data_8_8_0_sva_dfm_mx0;
  wire buf_acc_data_8_9_0_sva_dfm_mx0;
  wire buf_acc_data_8_10_0_sva_dfm_mx0;
  wire buf_acc_data_8_11_0_sva_dfm_mx0;
  wire buf_acc_data_8_12_0_sva_dfm_mx0;
  wire buf_acc_data_8_13_0_sva_dfm_mx0;
  wire buf_acc_data_8_14_0_sva_dfm_mx0;
  wire buf_acc_data_8_15_0_sva_dfm_mx0;
  wire buf_acc_data_8_16_0_sva_dfm_mx0;
  wire buf_acc_data_8_17_0_sva_dfm_mx0;
  wire buf_acc_data_9_0_0_sva_dfm_mx0;
  wire buf_acc_data_9_1_0_sva_dfm_mx0;
  wire buf_acc_data_9_2_0_sva_dfm_mx0;
  wire buf_acc_data_9_3_0_sva_dfm_mx0;
  wire buf_acc_data_9_4_0_sva_dfm_mx0;
  wire buf_acc_data_9_5_0_sva_dfm_mx0;
  wire buf_acc_data_9_6_0_sva_dfm_mx0;
  wire buf_acc_data_9_7_0_sva_dfm_mx0;
  wire buf_acc_data_9_8_0_sva_dfm_mx0;
  wire buf_acc_data_9_9_0_sva_dfm_mx0;
  wire buf_acc_data_9_10_0_sva_dfm_mx0;
  wire buf_acc_data_9_11_0_sva_dfm_mx0;
  wire buf_acc_data_9_12_0_sva_dfm_mx0;
  wire buf_acc_data_9_13_0_sva_dfm_mx0;
  wire buf_acc_data_9_14_0_sva_dfm_mx0;
  wire buf_acc_data_9_15_0_sva_dfm_mx0;
  wire buf_acc_data_9_16_0_sva_dfm_mx0;
  wire buf_acc_data_9_17_0_sva_dfm_mx0;
  wire buf_acc_data_10_0_0_sva_dfm_mx0;
  wire buf_acc_data_10_1_0_sva_dfm_mx0;
  wire buf_acc_data_10_2_0_sva_dfm_mx0;
  wire buf_acc_data_10_3_0_sva_dfm_mx0;
  wire buf_acc_data_10_4_0_sva_dfm_mx0;
  wire buf_acc_data_10_5_0_sva_dfm_mx0;
  wire buf_acc_data_10_6_0_sva_dfm_mx0;
  wire buf_acc_data_10_7_0_sva_dfm_mx0;
  wire buf_acc_data_10_8_0_sva_dfm_mx0;
  wire buf_acc_data_10_9_0_sva_dfm_mx0;
  wire buf_acc_data_10_10_0_sva_dfm_mx0;
  wire buf_acc_data_10_11_0_sva_dfm_mx0;
  wire buf_acc_data_10_12_0_sva_dfm_mx0;
  wire buf_acc_data_10_13_0_sva_dfm_mx0;
  wire buf_acc_data_10_14_0_sva_dfm_mx0;
  wire buf_acc_data_10_15_0_sva_dfm_mx0;
  wire buf_acc_data_10_16_0_sva_dfm_mx0;
  wire buf_acc_data_10_17_0_sva_dfm_mx0;
  wire buf_acc_data_11_0_0_sva_dfm_mx0;
  wire buf_acc_data_11_1_0_sva_dfm_mx0;
  wire buf_acc_data_11_2_0_sva_dfm_mx0;
  wire buf_acc_data_11_3_0_sva_dfm_mx0;
  wire buf_acc_data_11_4_0_sva_dfm_mx0;
  wire buf_acc_data_11_5_0_sva_dfm_mx0;
  wire buf_acc_data_11_6_0_sva_dfm_mx0;
  wire buf_acc_data_11_7_0_sva_dfm_mx0;
  wire buf_acc_data_11_8_0_sva_dfm_mx0;
  wire buf_acc_data_11_9_0_sva_dfm_mx0;
  wire buf_acc_data_11_10_0_sva_dfm_mx0;
  wire buf_acc_data_11_11_0_sva_dfm_mx0;
  wire buf_acc_data_11_12_0_sva_dfm_mx0;
  wire buf_acc_data_11_13_0_sva_dfm_mx0;
  wire buf_acc_data_11_14_0_sva_dfm_mx0;
  wire buf_acc_data_11_15_0_sva_dfm_mx0;
  wire buf_acc_data_11_16_0_sva_dfm_mx0;
  wire buf_acc_data_11_17_0_sva_dfm_mx0;
  wire buf_acc_data_12_0_0_sva_dfm_mx0;
  wire buf_acc_data_12_1_0_sva_dfm_mx0;
  wire buf_acc_data_12_2_0_sva_dfm_mx0;
  wire buf_acc_data_12_3_0_sva_dfm_mx0;
  wire buf_acc_data_12_4_0_sva_dfm_mx0;
  wire buf_acc_data_12_5_0_sva_dfm_mx0;
  wire buf_acc_data_12_6_0_sva_dfm_mx0;
  wire buf_acc_data_12_7_0_sva_dfm_mx0;
  wire buf_acc_data_12_8_0_sva_dfm_mx0;
  wire buf_acc_data_12_9_0_sva_dfm_mx0;
  wire buf_acc_data_12_10_0_sva_dfm_mx0;
  wire buf_acc_data_12_11_0_sva_dfm_mx0;
  wire buf_acc_data_12_12_0_sva_dfm_mx0;
  wire buf_acc_data_12_13_0_sva_dfm_mx0;
  wire buf_acc_data_12_14_0_sva_dfm_mx0;
  wire buf_acc_data_12_15_0_sva_dfm_mx0;
  wire buf_acc_data_12_16_0_sva_dfm_mx0;
  wire buf_acc_data_12_17_0_sva_dfm_mx0;
  wire buf_acc_data_13_0_0_sva_dfm_mx0;
  wire buf_acc_data_13_1_0_sva_dfm_mx0;
  wire buf_acc_data_13_2_0_sva_dfm_mx0;
  wire buf_acc_data_13_3_0_sva_dfm_mx0;
  wire buf_acc_data_13_4_0_sva_dfm_mx0;
  wire buf_acc_data_13_5_0_sva_dfm_mx0;
  wire buf_acc_data_13_6_0_sva_dfm_mx0;
  wire buf_acc_data_13_7_0_sva_dfm_mx0;
  wire buf_acc_data_13_8_0_sva_dfm_mx0;
  wire buf_acc_data_13_9_0_sva_dfm_mx0;
  wire buf_acc_data_13_10_0_sva_dfm_mx0;
  wire buf_acc_data_13_11_0_sva_dfm_mx0;
  wire buf_acc_data_13_12_0_sva_dfm_mx0;
  wire buf_acc_data_13_13_0_sva_dfm_mx0;
  wire buf_acc_data_13_14_0_sva_dfm_mx0;
  wire buf_acc_data_13_15_0_sva_dfm_mx0;
  wire buf_acc_data_13_16_0_sva_dfm_mx0;
  wire buf_acc_data_13_17_0_sva_dfm_mx0;
  wire buf_acc_data_14_0_0_sva_dfm_mx0;
  wire buf_acc_data_14_1_0_sva_dfm_mx0;
  wire buf_acc_data_14_2_0_sva_dfm_mx0;
  wire buf_acc_data_14_3_0_sva_dfm_mx0;
  wire buf_acc_data_14_4_0_sva_dfm_mx0;
  wire buf_acc_data_14_5_0_sva_dfm_mx0;
  wire buf_acc_data_14_6_0_sva_dfm_mx0;
  wire buf_acc_data_14_7_0_sva_dfm_mx0;
  wire buf_acc_data_14_8_0_sva_dfm_mx0;
  wire buf_acc_data_14_9_0_sva_dfm_mx0;
  wire buf_acc_data_14_10_0_sva_dfm_mx0;
  wire buf_acc_data_14_11_0_sva_dfm_mx0;
  wire buf_acc_data_14_12_0_sva_dfm_mx0;
  wire buf_acc_data_14_13_0_sva_dfm_mx0;
  wire buf_acc_data_14_14_0_sva_dfm_mx0;
  wire buf_acc_data_14_15_0_sva_dfm_mx0;
  wire buf_acc_data_14_16_0_sva_dfm_mx0;
  wire buf_acc_data_14_17_0_sva_dfm_mx0;
  wire buf_acc_data_15_0_0_sva_dfm_mx0;
  wire buf_acc_data_15_1_0_sva_dfm_mx0;
  wire buf_acc_data_15_2_0_sva_dfm_mx0;
  wire buf_acc_data_15_3_0_sva_dfm_mx0;
  wire buf_acc_data_15_4_0_sva_dfm_mx0;
  wire buf_acc_data_15_5_0_sva_dfm_mx0;
  wire buf_acc_data_15_6_0_sva_dfm_mx0;
  wire buf_acc_data_15_7_0_sva_dfm_mx0;
  wire buf_acc_data_15_8_0_sva_dfm_mx0;
  wire buf_acc_data_15_9_0_sva_dfm_mx0;
  wire buf_acc_data_15_10_0_sva_dfm_mx0;
  wire buf_acc_data_15_11_0_sva_dfm_mx0;
  wire buf_acc_data_15_12_0_sva_dfm_mx0;
  wire buf_acc_data_15_13_0_sva_dfm_mx0;
  wire buf_acc_data_15_14_0_sva_dfm_mx0;
  wire buf_acc_data_15_15_0_sva_dfm_mx0;
  wire buf_acc_data_15_16_0_sva_dfm_mx0;
  wire buf_acc_data_15_17_0_sva_dfm_mx0;
  wire buf_acc_data_16_0_0_sva_dfm_mx0;
  wire buf_acc_data_16_1_0_sva_dfm_mx0;
  wire buf_acc_data_16_2_0_sva_dfm_mx0;
  wire buf_acc_data_16_3_0_sva_dfm_mx0;
  wire buf_acc_data_16_4_0_sva_dfm_mx0;
  wire buf_acc_data_16_5_0_sva_dfm_mx0;
  wire buf_acc_data_16_6_0_sva_dfm_mx0;
  wire buf_acc_data_16_7_0_sva_dfm_mx0;
  wire buf_acc_data_16_8_0_sva_dfm_mx0;
  wire buf_acc_data_16_9_0_sva_dfm_mx0;
  wire buf_acc_data_16_10_0_sva_dfm_mx0;
  wire buf_acc_data_16_11_0_sva_dfm_mx0;
  wire buf_acc_data_16_12_0_sva_dfm_mx0;
  wire buf_acc_data_16_13_0_sva_dfm_mx0;
  wire buf_acc_data_16_14_0_sva_dfm_mx0;
  wire buf_acc_data_16_15_0_sva_dfm_mx0;
  wire buf_acc_data_16_16_0_sva_dfm_mx0;
  wire buf_acc_data_16_17_0_sva_dfm_mx0;
  wire buf_acc_data_17_0_0_sva_dfm_mx0;
  wire buf_acc_data_17_1_0_sva_dfm_mx0;
  wire buf_acc_data_17_2_0_sva_dfm_mx0;
  wire buf_acc_data_17_3_0_sva_dfm_mx0;
  wire buf_acc_data_17_4_0_sva_dfm_mx0;
  wire buf_acc_data_17_5_0_sva_dfm_mx0;
  wire buf_acc_data_17_6_0_sva_dfm_mx0;
  wire buf_acc_data_17_7_0_sva_dfm_mx0;
  wire buf_acc_data_17_8_0_sva_dfm_mx0;
  wire buf_acc_data_17_9_0_sva_dfm_mx0;
  wire buf_acc_data_17_10_0_sva_dfm_mx0;
  wire buf_acc_data_17_11_0_sva_dfm_mx0;
  wire buf_acc_data_17_12_0_sva_dfm_mx0;
  wire buf_acc_data_17_13_0_sva_dfm_mx0;
  wire buf_acc_data_17_14_0_sva_dfm_mx0;
  wire buf_acc_data_17_15_0_sva_dfm_mx0;
  wire buf_acc_data_17_16_0_sva_dfm_mx0;
  wire buf_acc_data_17_17_0_sva_dfm_mx0;
  wire [44:0] buf_acc_data_0_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_0_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_1_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_2_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_3_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_4_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_5_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_6_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_7_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_8_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_9_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_10_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_11_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_12_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_13_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_14_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_15_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_16_17_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_0_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_1_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_2_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_3_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_4_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_5_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_6_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_7_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_8_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_9_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_10_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_11_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_12_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_13_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_14_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_15_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_16_45_1_sva_dfm_1;
  wire [44:0] buf_acc_data_17_17_45_1_sva_dfm_1;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1;
  wire [4:0] PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5;
  wire [4:0] PADDING_LOOP_for_row_4_0_sva_2;
  wire [5:0] nl_PADDING_LOOP_for_row_4_0_sva_2;
  wire [4:0] PADDING_LOOP_for_for_col_4_0_sva_2;
  wire [5:0] nl_PADDING_LOOP_for_for_col_4_0_sva_2;
  wire [4:0] CONVOLUTION_LOOP_for_for_i_4_0_sva_2;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2;
  wire [3:0] nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_4;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2;
  wire [3:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_5;
  wire [13:0] STORE_LOOP_i_13_0_sva_2;
  wire [14:0] nl_STORE_LOOP_i_13_0_sva_2;
  wire STORE_LOOP_and_34_ssc_1;
  wire BATCH_LOOP_BATCH_LOOP_or_1_cse_1;
  wire BATCH_LOOP_BATCH_LOOP_or_2_cse_1;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_mx0;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_mx0;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1;
  wire [12:0] nl_CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_5_tmp_1;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_3;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1;
  wire CONVOLUTION_LOOP_for_for_for_asn_3570;
  wire CONVOLUTION_LOOP_for_for_for_asn_3572;
  wire CONVOLUTION_LOOP_for_for_for_asn_3574;
  wire CONVOLUTION_LOOP_for_for_for_asn_3576;
  wire CONVOLUTION_LOOP_for_for_for_asn_3578;
  wire CONVOLUTION_LOOP_for_for_for_asn_3580;
  wire CONVOLUTION_LOOP_for_for_for_asn_3582;
  wire CONVOLUTION_LOOP_for_for_for_asn_3584;
  wire CONVOLUTION_LOOP_for_for_for_asn_3586;
  wire CONVOLUTION_LOOP_for_for_for_asn_3588;
  wire CONVOLUTION_LOOP_for_for_for_asn_3590;
  wire CONVOLUTION_LOOP_for_for_for_asn_3592;
  wire CONVOLUTION_LOOP_for_for_for_asn_3594;
  wire CONVOLUTION_LOOP_for_for_for_asn_3596;
  wire CONVOLUTION_LOOP_for_for_for_asn_3598;
  wire CONVOLUTION_LOOP_for_for_for_asn_3600;
  wire CONVOLUTION_LOOP_for_for_for_asn_3602;
  wire CONVOLUTION_LOOP_for_for_for_asn_3604;
  wire CONVOLUTION_LOOP_for_for_for_asn_3606;
  wire CONVOLUTION_LOOP_for_for_for_asn_3608;
  wire CONVOLUTION_LOOP_for_for_for_asn_3610;
  wire CONVOLUTION_LOOP_for_for_for_asn_3612;
  wire CONVOLUTION_LOOP_for_for_for_asn_3614;
  wire CONVOLUTION_LOOP_for_for_for_asn_3616;
  wire CONVOLUTION_LOOP_for_for_for_asn_3618;
  wire CONVOLUTION_LOOP_for_for_for_asn_3620;
  wire CONVOLUTION_LOOP_for_for_for_asn_3622;
  wire CONVOLUTION_LOOP_for_for_for_asn_3624;
  wire CONVOLUTION_LOOP_for_for_for_asn_3626;
  wire CONVOLUTION_LOOP_for_for_for_asn_3628;
  wire CONVOLUTION_LOOP_for_for_for_asn_3630;
  wire CONVOLUTION_LOOP_for_for_for_asn_3632;
  wire CONVOLUTION_LOOP_for_for_for_asn_3634;
  wire CONVOLUTION_LOOP_for_for_for_asn_3636;
  wire CONVOLUTION_LOOP_for_for_for_asn_3638;
  wire CONVOLUTION_LOOP_for_for_for_asn_3640;
  wire CONVOLUTION_LOOP_for_for_for_asn_3642;
  wire CONVOLUTION_LOOP_for_for_for_asn_3644;
  wire CONVOLUTION_LOOP_for_for_for_asn_3646;
  wire CONVOLUTION_LOOP_for_for_for_asn_3648;
  wire CONVOLUTION_LOOP_for_for_for_asn_3650;
  wire CONVOLUTION_LOOP_for_for_for_asn_3652;
  wire CONVOLUTION_LOOP_for_for_for_asn_3654;
  wire CONVOLUTION_LOOP_for_for_for_asn_3656;
  wire CONVOLUTION_LOOP_for_for_for_asn_3658;
  wire CONVOLUTION_LOOP_for_for_for_asn_3660;
  wire CONVOLUTION_LOOP_for_for_for_asn_3662;
  wire CONVOLUTION_LOOP_for_for_for_asn_3664;
  wire CONVOLUTION_LOOP_for_for_for_asn_3666;
  wire CONVOLUTION_LOOP_for_for_for_asn_3668;
  wire CONVOLUTION_LOOP_for_for_for_asn_3670;
  wire CONVOLUTION_LOOP_for_for_for_asn_3672;
  wire CONVOLUTION_LOOP_for_for_for_asn_3674;
  wire CONVOLUTION_LOOP_for_for_for_asn_3676;
  wire CONVOLUTION_LOOP_for_for_for_asn_3678;
  wire CONVOLUTION_LOOP_for_for_for_asn_3680;
  wire CONVOLUTION_LOOP_for_for_for_asn_3682;
  wire CONVOLUTION_LOOP_for_for_for_asn_3684;
  wire CONVOLUTION_LOOP_for_for_for_asn_3686;
  wire CONVOLUTION_LOOP_for_for_for_asn_3688;
  wire CONVOLUTION_LOOP_for_for_for_asn_3690;
  wire CONVOLUTION_LOOP_for_for_for_asn_3692;
  wire CONVOLUTION_LOOP_for_for_for_asn_3694;
  wire CONVOLUTION_LOOP_for_for_for_asn_3696;
  wire CONVOLUTION_LOOP_for_for_for_asn_3698;
  wire CONVOLUTION_LOOP_for_for_for_asn_3700;
  wire CONVOLUTION_LOOP_for_for_for_asn_3702;
  wire CONVOLUTION_LOOP_for_for_for_asn_3704;
  wire CONVOLUTION_LOOP_for_for_for_asn_3706;
  wire CONVOLUTION_LOOP_for_for_for_asn_3708;
  wire CONVOLUTION_LOOP_for_for_for_asn_3710;
  wire CONVOLUTION_LOOP_for_for_for_asn_3712;
  wire CONVOLUTION_LOOP_for_for_for_asn_3714;
  wire CONVOLUTION_LOOP_for_for_for_asn_3716;
  wire CONVOLUTION_LOOP_for_for_for_asn_3718;
  wire CONVOLUTION_LOOP_for_for_for_asn_3720;
  wire CONVOLUTION_LOOP_for_for_for_asn_3722;
  wire CONVOLUTION_LOOP_for_for_for_asn_3724;
  wire CONVOLUTION_LOOP_for_for_for_asn_3726;
  wire CONVOLUTION_LOOP_for_for_for_asn_3728;
  wire CONVOLUTION_LOOP_for_for_for_asn_3730;
  wire CONVOLUTION_LOOP_for_for_for_asn_3732;
  wire CONVOLUTION_LOOP_for_for_for_asn_3734;
  wire CONVOLUTION_LOOP_for_for_for_asn_3736;
  wire CONVOLUTION_LOOP_for_for_for_asn_3738;
  wire CONVOLUTION_LOOP_for_for_for_asn_3740;
  wire CONVOLUTION_LOOP_for_for_for_asn_3742;
  wire CONVOLUTION_LOOP_for_for_for_asn_3744;
  wire CONVOLUTION_LOOP_for_for_for_asn_3746;
  wire CONVOLUTION_LOOP_for_for_for_asn_3748;
  wire CONVOLUTION_LOOP_for_for_for_asn_3750;
  wire CONVOLUTION_LOOP_for_for_for_asn_3752;
  wire CONVOLUTION_LOOP_for_for_for_asn_3754;
  wire CONVOLUTION_LOOP_for_for_for_asn_3756;
  wire CONVOLUTION_LOOP_for_for_for_asn_3758;
  wire CONVOLUTION_LOOP_for_for_for_asn_3760;
  wire CONVOLUTION_LOOP_for_for_for_asn_3762;
  wire CONVOLUTION_LOOP_for_for_for_asn_3764;
  wire CONVOLUTION_LOOP_for_for_for_asn_3766;
  wire CONVOLUTION_LOOP_for_for_for_asn_3768;
  wire CONVOLUTION_LOOP_for_for_for_asn_3770;
  wire CONVOLUTION_LOOP_for_for_for_asn_3772;
  wire CONVOLUTION_LOOP_for_for_for_asn_3774;
  wire CONVOLUTION_LOOP_for_for_for_asn_3776;
  wire CONVOLUTION_LOOP_for_for_for_asn_3778;
  wire CONVOLUTION_LOOP_for_for_for_asn_3780;
  wire CONVOLUTION_LOOP_for_for_for_asn_3782;
  wire CONVOLUTION_LOOP_for_for_for_asn_3784;
  wire CONVOLUTION_LOOP_for_for_for_asn_3786;
  wire CONVOLUTION_LOOP_for_for_for_asn_3788;
  wire CONVOLUTION_LOOP_for_for_for_asn_3790;
  wire CONVOLUTION_LOOP_for_for_for_asn_3792;
  wire CONVOLUTION_LOOP_for_for_for_asn_3794;
  wire CONVOLUTION_LOOP_for_for_for_asn_3796;
  wire CONVOLUTION_LOOP_for_for_for_asn_3798;
  wire CONVOLUTION_LOOP_for_for_for_asn_3800;
  wire CONVOLUTION_LOOP_for_for_for_asn_3802;
  wire CONVOLUTION_LOOP_for_for_for_asn_3804;
  wire CONVOLUTION_LOOP_for_for_for_asn_3806;
  wire CONVOLUTION_LOOP_for_for_for_asn_3808;
  wire CONVOLUTION_LOOP_for_for_for_asn_3810;
  wire CONVOLUTION_LOOP_for_for_for_asn_3812;
  wire CONVOLUTION_LOOP_for_for_for_asn_3814;
  wire CONVOLUTION_LOOP_for_for_for_asn_3816;
  wire CONVOLUTION_LOOP_for_for_for_asn_3818;
  wire CONVOLUTION_LOOP_for_for_for_asn_3820;
  wire CONVOLUTION_LOOP_for_for_for_asn_3822;
  wire CONVOLUTION_LOOP_for_for_for_asn_3824;
  wire CONVOLUTION_LOOP_for_for_for_asn_3826;
  wire CONVOLUTION_LOOP_for_for_for_asn_3828;
  wire CONVOLUTION_LOOP_for_for_for_asn_3830;
  wire CONVOLUTION_LOOP_for_for_for_asn_3832;
  wire CONVOLUTION_LOOP_for_for_for_asn_3834;
  wire CONVOLUTION_LOOP_for_for_for_asn_3836;
  wire CONVOLUTION_LOOP_for_for_for_asn_3838;
  wire CONVOLUTION_LOOP_for_for_for_asn_3840;
  wire CONVOLUTION_LOOP_for_for_for_asn_3842;
  wire CONVOLUTION_LOOP_for_for_for_asn_3844;
  wire CONVOLUTION_LOOP_for_for_for_asn_3846;
  wire CONVOLUTION_LOOP_for_for_for_asn_3848;
  wire CONVOLUTION_LOOP_for_for_for_asn_3850;
  wire CONVOLUTION_LOOP_for_for_for_asn_3852;
  wire CONVOLUTION_LOOP_for_for_for_asn_3854;
  wire CONVOLUTION_LOOP_for_for_for_asn_3856;
  wire CONVOLUTION_LOOP_for_for_for_asn_3858;
  wire CONVOLUTION_LOOP_for_for_for_asn_3860;
  wire CONVOLUTION_LOOP_for_for_for_asn_3862;
  wire CONVOLUTION_LOOP_for_for_for_asn_3864;
  wire CONVOLUTION_LOOP_for_for_for_asn_3866;
  wire CONVOLUTION_LOOP_for_for_for_asn_3868;
  wire CONVOLUTION_LOOP_for_for_for_asn_3870;
  wire CONVOLUTION_LOOP_for_for_for_asn_3872;
  wire CONVOLUTION_LOOP_for_for_for_asn_3874;
  wire CONVOLUTION_LOOP_for_for_for_asn_3876;
  wire CONVOLUTION_LOOP_for_for_for_asn_3878;
  wire CONVOLUTION_LOOP_for_for_for_asn_3880;
  wire CONVOLUTION_LOOP_for_for_for_asn_3882;
  wire CONVOLUTION_LOOP_for_for_for_asn_3884;
  wire CONVOLUTION_LOOP_for_for_for_asn_3886;
  wire CONVOLUTION_LOOP_for_for_for_asn_3888;
  wire CONVOLUTION_LOOP_for_for_for_asn_3890;
  wire CONVOLUTION_LOOP_for_for_for_asn_3892;
  wire CONVOLUTION_LOOP_for_for_for_asn_3894;
  wire CONVOLUTION_LOOP_for_for_for_asn_3896;
  wire CONVOLUTION_LOOP_for_for_for_asn_3898;
  wire CONVOLUTION_LOOP_for_for_for_asn_3900;
  wire CONVOLUTION_LOOP_for_for_for_asn_3902;
  wire CONVOLUTION_LOOP_for_for_for_asn_3904;
  wire CONVOLUTION_LOOP_for_for_for_asn_3906;
  wire CONVOLUTION_LOOP_for_for_for_asn_3908;
  wire CONVOLUTION_LOOP_for_for_for_asn_3910;
  wire CONVOLUTION_LOOP_for_for_for_asn_3912;
  wire CONVOLUTION_LOOP_for_for_for_asn_3914;
  wire CONVOLUTION_LOOP_for_for_for_asn_3916;
  wire CONVOLUTION_LOOP_for_for_for_asn_3918;
  wire CONVOLUTION_LOOP_for_for_for_asn_3920;
  wire CONVOLUTION_LOOP_for_for_for_asn_3922;
  wire CONVOLUTION_LOOP_for_for_for_asn_3924;
  wire CONVOLUTION_LOOP_for_for_for_asn_3926;
  wire CONVOLUTION_LOOP_for_for_for_asn_3928;
  wire CONVOLUTION_LOOP_for_for_for_asn_3930;
  wire CONVOLUTION_LOOP_for_for_for_asn_3932;
  wire CONVOLUTION_LOOP_for_for_for_asn_3934;
  wire CONVOLUTION_LOOP_for_for_for_asn_3936;
  wire CONVOLUTION_LOOP_for_for_for_asn_3938;
  wire CONVOLUTION_LOOP_for_for_for_asn_3940;
  wire CONVOLUTION_LOOP_for_for_for_asn_3942;
  wire CONVOLUTION_LOOP_for_for_for_asn_3944;
  wire CONVOLUTION_LOOP_for_for_for_asn_3946;
  wire CONVOLUTION_LOOP_for_for_for_asn_3948;
  wire CONVOLUTION_LOOP_for_for_for_asn_3950;
  wire CONVOLUTION_LOOP_for_for_for_asn_3952;
  wire CONVOLUTION_LOOP_for_for_for_asn_3954;
  wire CONVOLUTION_LOOP_for_for_for_asn_3956;
  wire CONVOLUTION_LOOP_for_for_for_asn_3958;
  wire CONVOLUTION_LOOP_for_for_for_asn_3960;
  wire CONVOLUTION_LOOP_for_for_for_asn_3962;
  wire CONVOLUTION_LOOP_for_for_for_asn_3964;
  wire CONVOLUTION_LOOP_for_for_for_asn_3966;
  wire CONVOLUTION_LOOP_for_for_for_asn_3968;
  wire CONVOLUTION_LOOP_for_for_for_asn_3970;
  wire CONVOLUTION_LOOP_for_for_for_asn_3972;
  wire CONVOLUTION_LOOP_for_for_for_asn_3974;
  wire CONVOLUTION_LOOP_for_for_for_asn_3976;
  wire CONVOLUTION_LOOP_for_for_for_asn_3978;
  wire CONVOLUTION_LOOP_for_for_for_asn_3980;
  wire CONVOLUTION_LOOP_for_for_for_asn_3982;
  wire CONVOLUTION_LOOP_for_for_for_asn_3984;
  wire CONVOLUTION_LOOP_for_for_for_asn_3986;
  wire CONVOLUTION_LOOP_for_for_for_asn_3988;
  wire CONVOLUTION_LOOP_for_for_for_asn_3990;
  wire CONVOLUTION_LOOP_for_for_for_asn_3992;
  wire CONVOLUTION_LOOP_for_for_for_asn_3994;
  wire CONVOLUTION_LOOP_for_for_for_asn_3996;
  wire CONVOLUTION_LOOP_for_for_for_asn_3998;
  wire CONVOLUTION_LOOP_for_for_for_asn_4000;
  wire CONVOLUTION_LOOP_for_for_for_asn_4002;
  wire CONVOLUTION_LOOP_for_for_for_asn_4004;
  wire CONVOLUTION_LOOP_for_for_for_asn_4006;
  wire CONVOLUTION_LOOP_for_for_for_asn_4008;
  wire CONVOLUTION_LOOP_for_for_for_asn_4010;
  wire CONVOLUTION_LOOP_for_for_for_asn_4012;
  wire CONVOLUTION_LOOP_for_for_for_asn_4014;
  wire CONVOLUTION_LOOP_for_for_for_asn_4016;
  wire CONVOLUTION_LOOP_for_for_for_asn_4018;
  wire CONVOLUTION_LOOP_for_for_for_asn_4020;
  wire CONVOLUTION_LOOP_for_for_for_asn_4022;
  wire CONVOLUTION_LOOP_for_for_for_asn_4024;
  wire CONVOLUTION_LOOP_for_for_for_asn_4026;
  wire CONVOLUTION_LOOP_for_for_for_asn_4028;
  wire CONVOLUTION_LOOP_for_for_for_asn_4030;
  wire CONVOLUTION_LOOP_for_for_for_asn_4032;
  wire CONVOLUTION_LOOP_for_for_for_asn_4034;
  wire CONVOLUTION_LOOP_for_for_for_asn_4036;
  wire CONVOLUTION_LOOP_for_for_for_asn_4038;
  wire CONVOLUTION_LOOP_for_for_for_asn_4040;
  wire CONVOLUTION_LOOP_for_for_for_asn_4042;
  wire CONVOLUTION_LOOP_for_for_for_asn_4044;
  wire CONVOLUTION_LOOP_for_for_for_asn_4046;
  wire CONVOLUTION_LOOP_for_for_for_asn_4048;
  wire CONVOLUTION_LOOP_for_for_for_asn_4050;
  wire CONVOLUTION_LOOP_for_for_for_asn_4052;
  wire CONVOLUTION_LOOP_for_for_for_asn_4054;
  wire CONVOLUTION_LOOP_for_for_for_asn_4056;
  wire CONVOLUTION_LOOP_for_for_for_asn_4058;
  wire CONVOLUTION_LOOP_for_for_for_asn_4060;
  wire CONVOLUTION_LOOP_for_for_for_asn_4062;
  wire CONVOLUTION_LOOP_for_for_for_asn_4064;
  wire CONVOLUTION_LOOP_for_for_for_asn_4066;
  wire CONVOLUTION_LOOP_for_for_for_asn_4068;
  wire CONVOLUTION_LOOP_for_for_for_asn_4070;
  wire CONVOLUTION_LOOP_for_for_for_asn_4072;
  wire CONVOLUTION_LOOP_for_for_for_asn_4074;
  wire CONVOLUTION_LOOP_for_for_for_asn_4076;
  wire CONVOLUTION_LOOP_for_for_for_asn_4078;
  wire CONVOLUTION_LOOP_for_for_for_asn_4080;
  wire CONVOLUTION_LOOP_for_for_for_asn_4082;
  wire CONVOLUTION_LOOP_for_for_for_asn_4084;
  wire CONVOLUTION_LOOP_for_for_for_asn_4086;
  wire CONVOLUTION_LOOP_for_for_for_asn_4088;
  wire CONVOLUTION_LOOP_for_for_for_asn_4090;
  wire CONVOLUTION_LOOP_for_for_for_asn_4092;
  wire CONVOLUTION_LOOP_for_for_for_asn_4094;
  wire CONVOLUTION_LOOP_for_for_for_asn_4096;
  wire CONVOLUTION_LOOP_for_for_for_asn_4098;
  wire CONVOLUTION_LOOP_for_for_for_asn_4100;
  wire CONVOLUTION_LOOP_for_for_for_asn_4102;
  wire CONVOLUTION_LOOP_for_for_for_asn_4104;
  wire CONVOLUTION_LOOP_for_for_for_asn_4106;
  wire CONVOLUTION_LOOP_for_for_for_asn_4108;
  wire CONVOLUTION_LOOP_for_for_for_asn_4110;
  wire CONVOLUTION_LOOP_for_for_for_asn_4112;
  wire CONVOLUTION_LOOP_for_for_for_asn_4114;
  wire CONVOLUTION_LOOP_for_for_for_asn_4116;
  wire CONVOLUTION_LOOP_for_for_for_asn_4118;
  wire CONVOLUTION_LOOP_for_for_for_asn_4120;
  wire CONVOLUTION_LOOP_for_for_for_asn_4122;
  wire CONVOLUTION_LOOP_for_for_for_asn_4124;
  wire CONVOLUTION_LOOP_for_for_for_asn_4126;
  wire CONVOLUTION_LOOP_for_for_for_asn_4128;
  wire CONVOLUTION_LOOP_for_for_for_asn_4130;
  wire CONVOLUTION_LOOP_for_for_for_asn_4132;
  wire CONVOLUTION_LOOP_for_for_for_asn_4134;
  wire CONVOLUTION_LOOP_for_for_for_asn_4136;
  wire CONVOLUTION_LOOP_for_for_for_asn_4138;
  wire CONVOLUTION_LOOP_for_for_for_asn_4140;
  wire CONVOLUTION_LOOP_for_for_for_asn_4142;
  wire CONVOLUTION_LOOP_for_for_for_asn_4144;
  wire CONVOLUTION_LOOP_for_for_for_asn_4146;
  wire CONVOLUTION_LOOP_for_for_for_asn_4148;
  wire CONVOLUTION_LOOP_for_for_for_asn_4150;
  wire CONVOLUTION_LOOP_for_for_for_asn_4152;
  wire CONVOLUTION_LOOP_for_for_for_asn_4154;
  wire CONVOLUTION_LOOP_for_for_for_asn_4156;
  wire CONVOLUTION_LOOP_for_for_for_asn_4158;
  wire CONVOLUTION_LOOP_for_for_for_asn_4160;
  wire CONVOLUTION_LOOP_for_for_for_asn_4162;
  wire CONVOLUTION_LOOP_for_for_for_asn_4164;
  wire CONVOLUTION_LOOP_for_for_for_asn_4166;
  wire CONVOLUTION_LOOP_for_for_for_asn_4168;
  wire CONVOLUTION_LOOP_for_for_for_asn_4170;
  wire CONVOLUTION_LOOP_for_for_for_asn_4172;
  wire CONVOLUTION_LOOP_for_for_for_asn_4174;
  wire CONVOLUTION_LOOP_for_for_for_asn_4176;
  wire CONVOLUTION_LOOP_for_for_for_asn_4178;
  wire CONVOLUTION_LOOP_for_for_for_asn_4180;
  wire CONVOLUTION_LOOP_for_for_for_asn_4182;
  wire CONVOLUTION_LOOP_for_for_for_asn_4184;
  wire CONVOLUTION_LOOP_for_for_for_asn_4186;
  wire CONVOLUTION_LOOP_for_for_for_asn_4188;
  wire CONVOLUTION_LOOP_for_for_for_asn_4190;
  wire CONVOLUTION_LOOP_for_for_for_asn_4192;
  wire CONVOLUTION_LOOP_for_for_for_asn_4194;
  wire CONVOLUTION_LOOP_for_for_for_asn_4196;
  wire CONVOLUTION_LOOP_for_for_for_asn_4198;
  wire CONVOLUTION_LOOP_for_for_for_asn_4200;
  wire CONVOLUTION_LOOP_for_for_for_asn_4202;
  wire CONVOLUTION_LOOP_for_for_for_asn_4204;
  wire CONVOLUTION_LOOP_for_for_for_asn_4206;
  wire CONVOLUTION_LOOP_for_for_for_asn_4208;
  wire CONVOLUTION_LOOP_for_for_for_asn_4210;
  wire CONVOLUTION_LOOP_for_for_for_asn_4212;
  wire CONVOLUTION_LOOP_for_for_for_asn_4214;
  wire CONVOLUTION_LOOP_for_for_for_asn_4216;
  wire CONVOLUTION_LOOP_for_for_for_asn_4218;
  wire CONVOLUTION_LOOP_for_for_for_asn_4220;
  wire CONVOLUTION_LOOP_for_for_for_asn_4222;
  wire CONVOLUTION_LOOP_for_for_for_asn_4224;
  wire CONVOLUTION_LOOP_for_for_for_asn_4226;
  wire CONVOLUTION_LOOP_for_for_for_asn_4228;
  wire CONVOLUTION_LOOP_for_for_for_asn_4230;
  wire CONVOLUTION_LOOP_for_for_for_asn_4232;
  wire CONVOLUTION_LOOP_for_for_for_asn_4234;
  wire CONVOLUTION_LOOP_for_for_for_asn_4236;
  wire CONVOLUTION_LOOP_for_for_for_asn_4238;
  wire CONVOLUTION_LOOP_for_for_for_asn_4240;
  wire CONVOLUTION_LOOP_for_for_for_asn_4242;
  wire CONVOLUTION_LOOP_for_for_for_asn_4244;
  wire CONVOLUTION_LOOP_for_for_for_asn_4246;
  wire CONVOLUTION_LOOP_for_for_for_asn_4248;
  wire CONVOLUTION_LOOP_for_for_for_asn_4250;
  wire CONVOLUTION_LOOP_for_for_for_asn_4252;
  wire CONVOLUTION_LOOP_for_for_for_asn_4254;
  wire CONVOLUTION_LOOP_for_for_for_asn_4256;
  wire CONVOLUTION_LOOP_for_for_for_asn_4258;
  wire CONVOLUTION_LOOP_for_for_for_asn_4260;
  wire CONVOLUTION_LOOP_for_for_for_asn_4262;
  wire CONVOLUTION_LOOP_for_for_for_asn_4264;
  wire CONVOLUTION_LOOP_for_for_for_asn_4266;
  wire CONVOLUTION_LOOP_for_for_for_asn_4268;
  wire CONVOLUTION_LOOP_for_for_for_asn_4270;
  wire CONVOLUTION_LOOP_for_for_for_asn_4272;
  wire CONVOLUTION_LOOP_for_for_for_asn_4274;
  wire CONVOLUTION_LOOP_for_for_for_asn_4276;
  wire CONVOLUTION_LOOP_for_for_for_asn_4278;
  wire CONVOLUTION_LOOP_for_for_for_asn_4280;
  wire CONVOLUTION_LOOP_for_for_for_asn_4282;
  wire CONVOLUTION_LOOP_for_for_for_asn_4284;
  wire CONVOLUTION_LOOP_for_for_for_asn_4286;
  wire CONVOLUTION_LOOP_for_for_for_asn_4288;
  wire CONVOLUTION_LOOP_for_for_for_asn_4290;
  wire CONVOLUTION_LOOP_for_for_for_asn_4292;
  wire CONVOLUTION_LOOP_for_for_for_asn_4294;
  wire CONVOLUTION_LOOP_for_for_for_asn_4296;
  wire CONVOLUTION_LOOP_for_for_for_asn_4298;
  wire CONVOLUTION_LOOP_for_for_for_asn_4300;
  wire CONVOLUTION_LOOP_for_for_for_asn_4302;
  wire CONVOLUTION_LOOP_for_for_for_asn_4304;
  wire CONVOLUTION_LOOP_for_for_for_asn_4306;
  wire CONVOLUTION_LOOP_for_for_for_asn_4308;
  wire CONVOLUTION_LOOP_for_for_for_asn_4310;
  wire CONVOLUTION_LOOP_for_for_for_asn_4312;
  wire CONVOLUTION_LOOP_for_for_for_asn_4314;
  wire CONVOLUTION_LOOP_for_for_for_asn_4316;
  wire CONVOLUTION_LOOP_for_for_for_asn_4318;
  wire CONVOLUTION_LOOP_for_for_for_asn_4320;
  wire CONVOLUTION_LOOP_for_for_for_asn_4322;
  wire CONVOLUTION_LOOP_for_for_for_asn_4324;
  wire CONVOLUTION_LOOP_for_for_for_asn_4326;
  wire CONVOLUTION_LOOP_for_for_for_asn_4328;
  wire CONVOLUTION_LOOP_for_for_for_asn_4330;
  wire CONVOLUTION_LOOP_for_for_for_asn_4332;
  wire CONVOLUTION_LOOP_for_for_for_asn_4334;
  wire CONVOLUTION_LOOP_for_for_for_asn_4336;
  wire CONVOLUTION_LOOP_for_for_for_asn_4338;
  wire CONVOLUTION_LOOP_for_for_for_asn_4340;
  wire CONVOLUTION_LOOP_for_for_for_asn_4342;
  wire CONVOLUTION_LOOP_for_for_for_asn_4344;
  wire CONVOLUTION_LOOP_for_for_for_asn_4346;
  wire CONVOLUTION_LOOP_for_for_for_asn_4348;
  wire CONVOLUTION_LOOP_for_for_for_asn_4350;
  wire CONVOLUTION_LOOP_for_for_for_asn_4352;
  wire CONVOLUTION_LOOP_for_for_for_asn_4354;
  wire CONVOLUTION_LOOP_for_for_for_asn_4356;
  wire CONVOLUTION_LOOP_for_for_for_asn_4358;
  wire CONVOLUTION_LOOP_for_for_for_asn_4360;
  wire CONVOLUTION_LOOP_for_for_for_asn_4362;
  wire CONVOLUTION_LOOP_for_for_for_asn_4364;
  wire CONVOLUTION_LOOP_for_for_for_asn_4366;
  wire CONVOLUTION_LOOP_for_for_for_asn_4368;
  wire CONVOLUTION_LOOP_for_for_for_asn_4370;
  wire CONVOLUTION_LOOP_for_for_for_asn_4372;
  wire CONVOLUTION_LOOP_for_for_for_asn_4374;
  wire CONVOLUTION_LOOP_for_for_for_asn_4376;
  wire CONVOLUTION_LOOP_for_for_for_asn_4378;
  wire CONVOLUTION_LOOP_for_for_for_asn_4380;
  wire CONVOLUTION_LOOP_for_for_for_asn_4382;
  wire CONVOLUTION_LOOP_for_for_for_asn_4384;
  wire CONVOLUTION_LOOP_for_for_for_asn_4386;
  wire CONVOLUTION_LOOP_for_for_for_asn_4388;
  wire CONVOLUTION_LOOP_for_for_for_asn_4390;
  wire CONVOLUTION_LOOP_for_for_for_asn_4392;
  wire CONVOLUTION_LOOP_for_for_for_asn_4394;
  wire CONVOLUTION_LOOP_for_for_for_asn_4396;
  wire CONVOLUTION_LOOP_for_for_for_asn_4398;
  wire CONVOLUTION_LOOP_for_for_for_asn_4400;
  wire CONVOLUTION_LOOP_for_for_for_asn_4402;
  wire CONVOLUTION_LOOP_for_for_for_asn_4404;
  wire CONVOLUTION_LOOP_for_for_for_asn_4406;
  wire CONVOLUTION_LOOP_for_for_for_asn_4408;
  wire CONVOLUTION_LOOP_for_for_for_asn_4410;
  wire CONVOLUTION_LOOP_for_for_for_asn_4412;
  wire CONVOLUTION_LOOP_for_for_for_asn_4414;
  wire CONVOLUTION_LOOP_for_for_for_asn_4416;
  wire CONVOLUTION_LOOP_for_for_for_asn_4418;
  wire CONVOLUTION_LOOP_for_for_for_asn_4420;
  wire CONVOLUTION_LOOP_for_for_for_asn_4422;
  wire CONVOLUTION_LOOP_for_for_for_asn_4424;
  wire CONVOLUTION_LOOP_for_for_for_asn_4426;
  wire CONVOLUTION_LOOP_for_for_for_asn_4428;
  wire CONVOLUTION_LOOP_for_for_for_asn_4430;
  wire CONVOLUTION_LOOP_for_for_for_asn_4432;
  wire CONVOLUTION_LOOP_for_for_for_asn_4434;
  wire CONVOLUTION_LOOP_for_for_for_asn_4436;
  wire CONVOLUTION_LOOP_for_for_for_asn_4438;
  wire CONVOLUTION_LOOP_for_for_for_asn_4440;
  wire CONVOLUTION_LOOP_for_for_for_asn_4442;
  wire CONVOLUTION_LOOP_for_for_for_asn_4444;
  wire CONVOLUTION_LOOP_for_for_for_asn_4446;
  wire CONVOLUTION_LOOP_for_for_for_asn_4448;
  wire CONVOLUTION_LOOP_for_for_for_asn_4450;
  wire CONVOLUTION_LOOP_for_for_for_asn_4452;
  wire CONVOLUTION_LOOP_for_for_for_asn_4454;
  wire CONVOLUTION_LOOP_for_for_for_asn_4456;
  wire CONVOLUTION_LOOP_for_for_for_asn_4458;
  wire CONVOLUTION_LOOP_for_for_for_asn_4460;
  wire CONVOLUTION_LOOP_for_for_for_asn_4462;
  wire CONVOLUTION_LOOP_for_for_for_asn_4464;
  wire CONVOLUTION_LOOP_for_for_for_asn_4466;
  wire CONVOLUTION_LOOP_for_for_for_asn_4468;
  wire CONVOLUTION_LOOP_for_for_for_asn_4470;
  wire CONVOLUTION_LOOP_for_for_for_asn_4472;
  wire CONVOLUTION_LOOP_for_for_for_asn_4474;
  wire CONVOLUTION_LOOP_for_for_for_asn_4476;
  wire CONVOLUTION_LOOP_for_for_for_asn_4478;
  wire CONVOLUTION_LOOP_for_for_for_asn_4480;
  wire CONVOLUTION_LOOP_for_for_for_asn_4482;
  wire CONVOLUTION_LOOP_for_for_for_asn_4484;
  wire CONVOLUTION_LOOP_for_for_for_asn_4486;
  wire CONVOLUTION_LOOP_for_for_for_asn_4488;
  wire CONVOLUTION_LOOP_for_for_for_asn_4490;
  wire CONVOLUTION_LOOP_for_for_for_asn_4492;
  wire CONVOLUTION_LOOP_for_for_for_asn_4494;
  wire CONVOLUTION_LOOP_for_for_for_asn_4496;
  wire CONVOLUTION_LOOP_for_for_for_asn_4498;
  wire CONVOLUTION_LOOP_for_for_for_asn_4500;
  wire CONVOLUTION_LOOP_for_for_for_asn_4502;
  wire CONVOLUTION_LOOP_for_for_for_asn_4504;
  wire CONVOLUTION_LOOP_for_for_for_asn_4506;
  wire CONVOLUTION_LOOP_for_for_for_asn_4508;
  wire CONVOLUTION_LOOP_for_for_for_asn_4510;
  wire CONVOLUTION_LOOP_for_for_for_asn_4512;
  wire CONVOLUTION_LOOP_for_for_for_asn_4514;
  wire CONVOLUTION_LOOP_for_for_for_asn_4516;
  wire CONVOLUTION_LOOP_for_for_for_asn_4518;
  wire CONVOLUTION_LOOP_for_for_for_asn_4520;
  wire CONVOLUTION_LOOP_for_for_for_asn_4522;
  wire CONVOLUTION_LOOP_for_for_for_asn_4524;
  wire CONVOLUTION_LOOP_for_for_for_asn_4526;
  wire CONVOLUTION_LOOP_for_for_for_asn_4528;
  wire CONVOLUTION_LOOP_for_for_for_asn_4530;
  wire CONVOLUTION_LOOP_for_for_for_asn_4532;
  wire CONVOLUTION_LOOP_for_for_for_asn_4534;
  wire CONVOLUTION_LOOP_for_for_for_asn_4536;
  wire CONVOLUTION_LOOP_for_for_for_asn_4538;
  wire CONVOLUTION_LOOP_for_for_for_asn_4540;
  wire CONVOLUTION_LOOP_for_for_for_asn_4542;
  wire CONVOLUTION_LOOP_for_for_for_asn_4544;
  wire CONVOLUTION_LOOP_for_for_for_asn_4546;
  wire CONVOLUTION_LOOP_for_for_for_asn_4548;
  wire CONVOLUTION_LOOP_for_for_for_asn_4550;
  wire CONVOLUTION_LOOP_for_for_for_asn_4552;
  wire CONVOLUTION_LOOP_for_for_for_asn_4554;
  wire CONVOLUTION_LOOP_for_for_for_asn_4556;
  wire CONVOLUTION_LOOP_for_for_for_asn_4558;
  wire CONVOLUTION_LOOP_for_for_for_asn_4560;
  wire CONVOLUTION_LOOP_for_for_for_asn_4562;
  wire CONVOLUTION_LOOP_for_for_for_asn_4564;
  wire CONVOLUTION_LOOP_for_for_for_asn_4566;
  wire CONVOLUTION_LOOP_for_for_for_asn_4568;
  wire CONVOLUTION_LOOP_for_for_for_asn_4570;
  wire CONVOLUTION_LOOP_for_for_for_asn_4572;
  wire CONVOLUTION_LOOP_for_for_for_asn_4574;
  wire CONVOLUTION_LOOP_for_for_for_asn_4576;
  wire CONVOLUTION_LOOP_for_for_for_asn_4578;
  wire CONVOLUTION_LOOP_for_for_for_asn_4580;
  wire CONVOLUTION_LOOP_for_for_for_asn_4582;
  wire CONVOLUTION_LOOP_for_for_for_asn_4584;
  wire CONVOLUTION_LOOP_for_for_for_asn_4586;
  wire CONVOLUTION_LOOP_for_for_for_asn_4588;
  wire CONVOLUTION_LOOP_for_for_for_asn_4590;
  wire CONVOLUTION_LOOP_for_for_for_asn_4592;
  wire CONVOLUTION_LOOP_for_for_for_asn_4594;
  wire CONVOLUTION_LOOP_for_for_for_asn_4596;
  wire CONVOLUTION_LOOP_for_for_for_asn_4598;
  wire CONVOLUTION_LOOP_for_for_for_asn_4600;
  wire CONVOLUTION_LOOP_for_for_for_asn_4602;
  wire CONVOLUTION_LOOP_for_for_for_asn_4604;
  wire CONVOLUTION_LOOP_for_for_for_asn_4606;
  wire CONVOLUTION_LOOP_for_for_for_asn_4608;
  wire CONVOLUTION_LOOP_for_for_for_asn_4610;
  wire CONVOLUTION_LOOP_for_for_for_asn_4612;
  wire CONVOLUTION_LOOP_for_for_for_asn_4614;
  wire CONVOLUTION_LOOP_for_for_for_asn_4616;
  wire CONVOLUTION_LOOP_for_for_for_asn_4618;
  wire CONVOLUTION_LOOP_for_for_for_asn_4620;
  wire CONVOLUTION_LOOP_for_for_for_asn_4622;
  wire CONVOLUTION_LOOP_for_for_for_asn_4624;
  wire CONVOLUTION_LOOP_for_for_for_asn_4626;
  wire CONVOLUTION_LOOP_for_for_for_asn_4628;
  wire CONVOLUTION_LOOP_for_for_for_asn_4630;
  wire CONVOLUTION_LOOP_for_for_for_asn_4632;
  wire CONVOLUTION_LOOP_for_for_for_asn_4634;
  wire CONVOLUTION_LOOP_for_for_for_asn_4636;
  wire CONVOLUTION_LOOP_for_for_for_asn_4638;
  wire CONVOLUTION_LOOP_for_for_for_asn_4640;
  wire CONVOLUTION_LOOP_for_for_for_asn_4642;
  wire CONVOLUTION_LOOP_for_for_for_asn_4644;
  wire CONVOLUTION_LOOP_for_for_for_asn_4646;
  wire CONVOLUTION_LOOP_for_for_for_asn_4648;
  wire CONVOLUTION_LOOP_for_for_for_asn_4650;
  wire CONVOLUTION_LOOP_for_for_for_asn_4652;
  wire CONVOLUTION_LOOP_for_for_for_asn_4654;
  wire CONVOLUTION_LOOP_for_for_for_asn_4656;
  wire CONVOLUTION_LOOP_for_for_for_asn_4658;
  wire CONVOLUTION_LOOP_for_for_for_asn_4660;
  wire CONVOLUTION_LOOP_for_for_for_asn_4662;
  wire CONVOLUTION_LOOP_for_for_for_asn_4664;
  wire CONVOLUTION_LOOP_for_for_for_asn_4666;
  wire CONVOLUTION_LOOP_for_for_for_asn_4668;
  wire CONVOLUTION_LOOP_for_for_for_asn_4670;
  wire CONVOLUTION_LOOP_for_for_for_asn_4672;
  wire CONVOLUTION_LOOP_for_for_for_asn_4674;
  wire CONVOLUTION_LOOP_for_for_for_asn_4676;
  wire CONVOLUTION_LOOP_for_for_for_asn_4678;
  wire CONVOLUTION_LOOP_for_for_for_asn_4680;
  wire CONVOLUTION_LOOP_for_for_for_asn_4682;
  wire CONVOLUTION_LOOP_for_for_for_asn_4684;
  wire CONVOLUTION_LOOP_for_for_for_asn_4686;
  wire CONVOLUTION_LOOP_for_for_for_asn_4688;
  wire CONVOLUTION_LOOP_for_for_for_asn_4690;
  wire CONVOLUTION_LOOP_for_for_for_asn_4692;
  wire CONVOLUTION_LOOP_for_for_for_asn_4694;
  wire CONVOLUTION_LOOP_for_for_for_asn_4696;
  wire CONVOLUTION_LOOP_for_for_for_asn_4698;
  wire CONVOLUTION_LOOP_for_for_for_asn_4700;
  wire CONVOLUTION_LOOP_for_for_for_asn_4702;
  wire CONVOLUTION_LOOP_for_for_for_asn_4704;
  wire CONVOLUTION_LOOP_for_for_for_asn_4706;
  wire CONVOLUTION_LOOP_for_for_for_asn_4708;
  wire CONVOLUTION_LOOP_for_for_for_asn_4710;
  wire CONVOLUTION_LOOP_for_for_for_asn_4712;
  wire CONVOLUTION_LOOP_for_for_for_asn_4714;
  wire CONVOLUTION_LOOP_for_for_for_asn_4716;
  wire CONVOLUTION_LOOP_for_for_for_asn_4718;
  wire CONVOLUTION_LOOP_for_for_for_asn_4720;
  wire CONVOLUTION_LOOP_for_for_for_asn_4722;
  wire CONVOLUTION_LOOP_for_for_for_asn_4724;
  wire CONVOLUTION_LOOP_for_for_for_asn_4726;
  wire CONVOLUTION_LOOP_for_for_for_asn_4728;
  wire CONVOLUTION_LOOP_for_for_for_asn_4730;
  wire CONVOLUTION_LOOP_for_for_for_asn_4732;
  wire CONVOLUTION_LOOP_for_for_for_asn_4734;
  wire CONVOLUTION_LOOP_for_for_for_asn_4736;
  wire CONVOLUTION_LOOP_for_for_for_asn_4738;
  wire CONVOLUTION_LOOP_for_for_for_asn_4740;
  wire CONVOLUTION_LOOP_for_for_for_asn_4742;
  wire CONVOLUTION_LOOP_for_for_for_asn_4744;
  wire CONVOLUTION_LOOP_for_for_for_asn_4746;
  wire CONVOLUTION_LOOP_for_for_for_asn_4748;
  wire CONVOLUTION_LOOP_for_for_for_asn_4750;
  wire CONVOLUTION_LOOP_for_for_for_asn_4752;
  wire CONVOLUTION_LOOP_for_for_for_asn_4754;
  wire CONVOLUTION_LOOP_for_for_for_asn_4756;
  wire CONVOLUTION_LOOP_for_for_for_asn_4758;
  wire CONVOLUTION_LOOP_for_for_for_asn_4760;
  wire CONVOLUTION_LOOP_for_for_for_asn_4762;
  wire CONVOLUTION_LOOP_for_for_for_asn_4764;
  wire CONVOLUTION_LOOP_for_for_for_asn_4766;
  wire CONVOLUTION_LOOP_for_for_for_asn_4768;
  wire CONVOLUTION_LOOP_for_for_for_asn_4770;
  wire CONVOLUTION_LOOP_for_for_for_asn_4772;
  wire CONVOLUTION_LOOP_for_for_for_asn_4774;
  wire CONVOLUTION_LOOP_for_for_for_asn_4776;
  wire CONVOLUTION_LOOP_for_for_for_asn_4778;
  wire CONVOLUTION_LOOP_for_for_for_asn_4780;
  wire CONVOLUTION_LOOP_for_for_for_asn_4782;
  wire CONVOLUTION_LOOP_for_for_for_asn_4784;
  wire CONVOLUTION_LOOP_for_for_for_asn_4786;
  wire CONVOLUTION_LOOP_for_for_for_asn_4788;
  wire CONVOLUTION_LOOP_for_for_for_asn_4790;
  wire CONVOLUTION_LOOP_for_for_for_asn_4792;
  wire CONVOLUTION_LOOP_for_for_for_asn_4794;
  wire CONVOLUTION_LOOP_for_for_for_asn_4796;
  wire CONVOLUTION_LOOP_for_for_for_asn_4798;
  wire CONVOLUTION_LOOP_for_for_for_asn_4800;
  wire CONVOLUTION_LOOP_for_for_for_asn_4802;
  wire CONVOLUTION_LOOP_for_for_for_asn_4804;
  wire CONVOLUTION_LOOP_for_for_for_asn_4806;
  wire CONVOLUTION_LOOP_for_for_for_asn_4808;
  wire CONVOLUTION_LOOP_for_for_for_asn_4810;
  wire CONVOLUTION_LOOP_for_for_for_asn_4812;
  wire CONVOLUTION_LOOP_for_for_for_asn_4814;
  wire CONVOLUTION_LOOP_for_for_for_asn_4816;
  wire CONVOLUTION_LOOP_for_for_for_asn_4818;
  wire CONVOLUTION_LOOP_for_for_for_asn_4820;
  wire CONVOLUTION_LOOP_for_for_for_asn_4822;
  wire CONVOLUTION_LOOP_for_for_for_asn_4824;
  wire CONVOLUTION_LOOP_for_for_for_asn_4826;
  wire CONVOLUTION_LOOP_for_for_for_asn_4828;
  wire CONVOLUTION_LOOP_for_for_for_asn_4830;
  wire CONVOLUTION_LOOP_for_for_for_asn_4832;
  wire CONVOLUTION_LOOP_for_for_for_asn_4834;
  wire CONVOLUTION_LOOP_for_for_for_asn_4836;
  wire CONVOLUTION_LOOP_for_for_for_asn_4838;
  wire CONVOLUTION_LOOP_for_for_for_asn_4840;
  wire CONVOLUTION_LOOP_for_for_for_asn_4842;
  wire CONVOLUTION_LOOP_for_for_for_asn_4844;
  wire CONVOLUTION_LOOP_for_for_for_asn_4846;
  wire CONVOLUTION_LOOP_for_for_for_asn_4848;
  wire CONVOLUTION_LOOP_for_for_for_asn_4850;
  wire CONVOLUTION_LOOP_for_for_for_asn_4852;
  wire CONVOLUTION_LOOP_for_for_for_asn_4854;
  wire CONVOLUTION_LOOP_for_for_for_asn_4856;
  wire CONVOLUTION_LOOP_for_for_for_asn_4858;
  wire CONVOLUTION_LOOP_for_for_for_asn_4860;
  wire CONVOLUTION_LOOP_for_for_for_asn_4862;
  wire CONVOLUTION_LOOP_for_for_for_asn_4864;
  wire CONVOLUTION_LOOP_for_for_for_asn_4866;
  wire CONVOLUTION_LOOP_for_for_for_asn_4868;
  wire CONVOLUTION_LOOP_for_for_for_asn_4870;
  wire CONVOLUTION_LOOP_for_for_for_asn_4872;
  wire CONVOLUTION_LOOP_for_for_for_asn_4874;
  wire CONVOLUTION_LOOP_for_for_for_asn_4876;
  wire CONVOLUTION_LOOP_for_for_for_asn_4878;
  wire CONVOLUTION_LOOP_for_for_for_asn_4880;
  wire CONVOLUTION_LOOP_for_for_for_asn_4882;
  wire CONVOLUTION_LOOP_for_for_for_asn_4884;
  wire CONVOLUTION_LOOP_for_for_for_asn_4886;
  wire CONVOLUTION_LOOP_for_for_for_asn_4888;
  wire CONVOLUTION_LOOP_for_for_for_asn_4890;
  wire CONVOLUTION_LOOP_for_for_for_asn_4892;
  wire CONVOLUTION_LOOP_for_for_for_asn_4894;
  wire CONVOLUTION_LOOP_for_for_for_asn_4896;
  wire CONVOLUTION_LOOP_for_for_for_asn_4898;
  wire CONVOLUTION_LOOP_for_for_for_asn_4900;
  wire CONVOLUTION_LOOP_for_for_for_asn_4902;
  wire CONVOLUTION_LOOP_for_for_for_asn_4904;
  wire CONVOLUTION_LOOP_for_for_for_asn_4906;
  wire CONVOLUTION_LOOP_for_for_for_asn_4908;
  wire CONVOLUTION_LOOP_for_for_for_asn_4910;
  wire CONVOLUTION_LOOP_for_for_for_asn_4912;
  wire CONVOLUTION_LOOP_for_for_for_asn_4914;
  wire CONVOLUTION_LOOP_for_for_for_asn_4916;
  wire CONVOLUTION_LOOP_for_for_for_asn_4918;
  wire CONVOLUTION_LOOP_for_for_for_asn_4920;
  wire CONVOLUTION_LOOP_for_for_for_asn_4922;
  wire CONVOLUTION_LOOP_for_for_for_asn_4924;
  wire CONVOLUTION_LOOP_for_for_for_asn_4926;
  wire CONVOLUTION_LOOP_for_for_for_asn_4928;
  wire CONVOLUTION_LOOP_for_for_for_asn_4930;
  wire CONVOLUTION_LOOP_for_for_for_asn_4932;
  wire CONVOLUTION_LOOP_for_for_for_asn_4934;
  wire CONVOLUTION_LOOP_for_for_for_asn_4936;
  wire CONVOLUTION_LOOP_for_for_for_asn_4938;
  wire CONVOLUTION_LOOP_for_for_for_asn_4940;
  wire CONVOLUTION_LOOP_for_for_for_asn_4942;
  wire CONVOLUTION_LOOP_for_for_for_asn_4944;
  wire CONVOLUTION_LOOP_for_for_for_asn_4946;
  wire CONVOLUTION_LOOP_for_for_for_asn_4948;
  wire CONVOLUTION_LOOP_for_for_for_asn_4950;
  wire CONVOLUTION_LOOP_for_for_for_asn_4952;
  wire CONVOLUTION_LOOP_for_for_for_asn_4954;
  wire CONVOLUTION_LOOP_for_for_for_asn_4956;
  wire CONVOLUTION_LOOP_for_for_for_asn_4958;
  wire CONVOLUTION_LOOP_for_for_for_asn_4960;
  wire CONVOLUTION_LOOP_for_for_for_asn_4962;
  wire CONVOLUTION_LOOP_for_for_for_asn_4964;
  wire CONVOLUTION_LOOP_for_for_for_asn_4966;
  wire CONVOLUTION_LOOP_for_for_for_asn_4968;
  wire CONVOLUTION_LOOP_for_for_for_asn_4970;
  wire CONVOLUTION_LOOP_for_for_for_asn_4972;
  wire CONVOLUTION_LOOP_for_for_for_asn_4974;
  wire CONVOLUTION_LOOP_for_for_for_asn_4976;
  wire CONVOLUTION_LOOP_for_for_for_asn_4978;
  wire CONVOLUTION_LOOP_for_for_for_asn_4980;
  wire CONVOLUTION_LOOP_for_for_for_asn_4982;
  wire CONVOLUTION_LOOP_for_for_for_asn_4984;
  wire CONVOLUTION_LOOP_for_for_for_asn_4986;
  wire CONVOLUTION_LOOP_for_for_for_asn_4988;
  wire CONVOLUTION_LOOP_for_for_for_asn_4990;
  wire CONVOLUTION_LOOP_for_for_for_asn_4992;
  wire CONVOLUTION_LOOP_for_for_for_asn_4994;
  wire CONVOLUTION_LOOP_for_for_for_asn_4996;
  wire CONVOLUTION_LOOP_for_for_for_asn_4998;
  wire CONVOLUTION_LOOP_for_for_for_asn_5000;
  wire CONVOLUTION_LOOP_for_for_for_asn_5002;
  wire CONVOLUTION_LOOP_for_for_for_asn_5004;
  wire CONVOLUTION_LOOP_for_for_for_asn_5006;
  wire CONVOLUTION_LOOP_for_for_for_asn_5008;
  wire CONVOLUTION_LOOP_for_for_for_asn_5010;
  wire CONVOLUTION_LOOP_for_for_for_asn_5012;
  wire CONVOLUTION_LOOP_for_for_for_asn_5014;
  wire CONVOLUTION_LOOP_for_for_for_asn_5016;
  wire CONVOLUTION_LOOP_for_for_for_asn_5018;
  wire CONVOLUTION_LOOP_for_for_for_asn_5020;
  wire CONVOLUTION_LOOP_for_for_for_asn_5022;
  wire CONVOLUTION_LOOP_for_for_for_asn_5024;
  wire CONVOLUTION_LOOP_for_for_for_asn_5026;
  wire CONVOLUTION_LOOP_for_for_for_asn_5028;
  wire CONVOLUTION_LOOP_for_for_for_asn_5030;
  wire CONVOLUTION_LOOP_for_for_for_asn_5032;
  wire CONVOLUTION_LOOP_for_for_for_asn_5034;
  wire CONVOLUTION_LOOP_for_for_for_asn_5036;
  wire CONVOLUTION_LOOP_for_for_for_asn_5038;
  wire CONVOLUTION_LOOP_for_for_for_asn_5040;
  wire CONVOLUTION_LOOP_for_for_for_asn_5042;
  wire CONVOLUTION_LOOP_for_for_for_asn_5044;
  wire CONVOLUTION_LOOP_for_for_for_asn_5046;
  wire CONVOLUTION_LOOP_for_for_for_asn_5048;
  wire CONVOLUTION_LOOP_for_for_for_asn_5050;
  wire CONVOLUTION_LOOP_for_for_for_asn_5052;
  wire CONVOLUTION_LOOP_for_for_for_asn_5054;
  wire CONVOLUTION_LOOP_for_for_for_asn_5056;
  wire CONVOLUTION_LOOP_for_for_for_asn_5058;
  wire CONVOLUTION_LOOP_for_for_for_asn_5060;
  wire CONVOLUTION_LOOP_for_for_for_asn_5062;
  wire CONVOLUTION_LOOP_for_for_for_asn_5064;
  wire CONVOLUTION_LOOP_for_for_for_asn_5066;
  wire CONVOLUTION_LOOP_for_for_for_asn_5068;
  wire CONVOLUTION_LOOP_for_for_for_asn_5070;
  wire CONVOLUTION_LOOP_for_for_for_asn_5072;
  wire CONVOLUTION_LOOP_for_for_for_asn_5074;
  wire CONVOLUTION_LOOP_for_for_for_asn_5076;
  wire CONVOLUTION_LOOP_for_for_for_asn_5078;
  wire CONVOLUTION_LOOP_for_for_for_asn_5080;
  wire CONVOLUTION_LOOP_for_for_for_asn_5082;
  wire CONVOLUTION_LOOP_for_for_for_asn_5084;
  wire CONVOLUTION_LOOP_for_for_for_asn_5086;
  wire CONVOLUTION_LOOP_for_for_for_asn_5088;
  wire CONVOLUTION_LOOP_for_for_for_asn_5090;
  wire CONVOLUTION_LOOP_for_for_for_asn_5092;
  wire CONVOLUTION_LOOP_for_for_for_asn_5094;
  wire CONVOLUTION_LOOP_for_for_for_asn_5096;
  wire CONVOLUTION_LOOP_for_for_for_asn_5098;
  wire CONVOLUTION_LOOP_for_for_for_asn_5100;
  wire CONVOLUTION_LOOP_for_for_for_asn_5102;
  wire CONVOLUTION_LOOP_for_for_for_asn_5104;
  wire CONVOLUTION_LOOP_for_for_for_asn_5106;
  wire CONVOLUTION_LOOP_for_for_for_asn_5108;
  wire CONVOLUTION_LOOP_for_for_for_asn_5110;
  wire CONVOLUTION_LOOP_for_for_for_asn_5112;
  wire CONVOLUTION_LOOP_for_for_for_asn_5114;
  wire CONVOLUTION_LOOP_for_for_for_asn_5116;
  wire CONVOLUTION_LOOP_for_for_for_asn_5118;
  wire CONVOLUTION_LOOP_for_for_for_asn_5120;
  wire CONVOLUTION_LOOP_for_for_for_asn_5122;
  wire CONVOLUTION_LOOP_for_for_for_asn_5124;
  wire CONVOLUTION_LOOP_for_for_for_asn_5126;
  wire CONVOLUTION_LOOP_for_for_for_asn_5128;
  wire CONVOLUTION_LOOP_for_for_for_asn_5130;
  wire CONVOLUTION_LOOP_for_for_for_asn_5132;
  wire CONVOLUTION_LOOP_for_for_for_asn_5134;
  wire CONVOLUTION_LOOP_for_for_for_asn_5136;
  wire CONVOLUTION_LOOP_for_for_for_asn_5138;
  wire CONVOLUTION_LOOP_for_for_for_asn_5140;
  wire CONVOLUTION_LOOP_for_for_for_asn_5142;
  wire CONVOLUTION_LOOP_for_for_for_asn_5144;
  wire CONVOLUTION_LOOP_for_for_for_asn_5146;
  wire CONVOLUTION_LOOP_for_for_for_asn_5148;
  wire CONVOLUTION_LOOP_for_for_for_asn_5150;
  wire CONVOLUTION_LOOP_for_for_for_asn_5152;
  wire CONVOLUTION_LOOP_for_for_for_asn_5154;
  wire CONVOLUTION_LOOP_for_for_for_asn_5156;
  wire CONVOLUTION_LOOP_for_for_for_asn_5158;
  wire CONVOLUTION_LOOP_for_for_for_asn_5160;
  wire CONVOLUTION_LOOP_for_for_for_asn_5162;
  wire CONVOLUTION_LOOP_for_for_for_asn_5164;
  wire CONVOLUTION_LOOP_for_for_for_asn_5166;
  wire CONVOLUTION_LOOP_for_for_for_asn_5168;
  wire CONVOLUTION_LOOP_for_for_for_asn_5170;
  wire CONVOLUTION_LOOP_for_for_for_asn_5172;
  wire CONVOLUTION_LOOP_for_for_for_asn_5174;
  wire CONVOLUTION_LOOP_for_for_for_asn_5176;
  wire CONVOLUTION_LOOP_for_for_for_asn_5178;
  wire CONVOLUTION_LOOP_for_for_for_asn_5180;
  wire CONVOLUTION_LOOP_for_for_for_asn_5182;
  wire CONVOLUTION_LOOP_for_for_for_asn_5184;
  wire CONVOLUTION_LOOP_for_for_for_asn_5186;
  wire CONVOLUTION_LOOP_for_for_for_asn_5188;
  wire CONVOLUTION_LOOP_for_for_for_asn_5190;
  wire CONVOLUTION_LOOP_for_for_for_asn_5192;
  wire CONVOLUTION_LOOP_for_for_for_asn_5194;
  wire CONVOLUTION_LOOP_for_for_for_asn_5196;
  wire CONVOLUTION_LOOP_for_for_for_asn_5198;
  wire CONVOLUTION_LOOP_for_for_for_asn_5200;
  wire CONVOLUTION_LOOP_for_for_for_asn_5202;
  wire CONVOLUTION_LOOP_for_for_for_asn_5204;
  wire CONVOLUTION_LOOP_for_for_for_asn_5206;
  wire CONVOLUTION_LOOP_for_for_for_asn_5208;
  wire CONVOLUTION_LOOP_for_for_for_asn_5210;
  wire CONVOLUTION_LOOP_for_for_for_asn_5212;
  wire CONVOLUTION_LOOP_for_for_for_asn_5214;
  wire CONVOLUTION_LOOP_for_for_for_asn_5216;
  wire CONVOLUTION_LOOP_for_for_for_asn_5218;
  wire CONVOLUTION_LOOP_for_for_for_asn_5220;
  wire CONVOLUTION_LOOP_for_for_for_asn_5222;
  wire CONVOLUTION_LOOP_for_for_for_asn_5224;
  wire CONVOLUTION_LOOP_for_for_for_asn_5226;
  wire CONVOLUTION_LOOP_for_for_for_asn_5228;
  wire CONVOLUTION_LOOP_for_for_for_asn_5230;
  wire CONVOLUTION_LOOP_for_for_for_asn_5232;
  wire CONVOLUTION_LOOP_for_for_for_asn_5234;
  wire CONVOLUTION_LOOP_for_for_for_asn_5236;
  wire CONVOLUTION_LOOP_for_for_for_asn_5238;
  wire CONVOLUTION_LOOP_for_for_for_asn_5240;
  wire CONVOLUTION_LOOP_for_for_for_asn_5242;
  wire CONVOLUTION_LOOP_for_for_for_asn_5244;
  wire CONVOLUTION_LOOP_for_for_for_asn_5246;
  wire CONVOLUTION_LOOP_for_for_for_asn_5248;
  wire CONVOLUTION_LOOP_for_for_for_asn_5250;
  wire CONVOLUTION_LOOP_for_for_for_asn_5252;
  wire CONVOLUTION_LOOP_for_for_for_asn_5254;
  wire CONVOLUTION_LOOP_for_for_for_asn_5256;
  wire CONVOLUTION_LOOP_for_for_for_asn_5258;
  wire CONVOLUTION_LOOP_for_for_for_asn_5260;
  wire CONVOLUTION_LOOP_for_for_for_asn_5262;
  wire CONVOLUTION_LOOP_for_for_for_asn_5264;
  wire CONVOLUTION_LOOP_for_for_for_asn_5266;
  wire CONVOLUTION_LOOP_for_for_for_asn_5268;
  wire CONVOLUTION_LOOP_for_for_for_asn_5270;
  wire CONVOLUTION_LOOP_for_for_for_asn_5272;
  wire CONVOLUTION_LOOP_for_for_for_asn_5274;
  wire CONVOLUTION_LOOP_for_for_for_asn_5276;
  wire CONVOLUTION_LOOP_for_for_for_asn_5278;
  wire CONVOLUTION_LOOP_for_for_for_asn_5280;
  wire CONVOLUTION_LOOP_for_for_for_asn_5282;
  wire CONVOLUTION_LOOP_for_for_for_asn_5284;
  wire CONVOLUTION_LOOP_for_for_for_asn_5286;
  wire CONVOLUTION_LOOP_for_for_for_asn_5288;
  wire CONVOLUTION_LOOP_for_for_for_asn_5290;
  wire CONVOLUTION_LOOP_for_for_for_asn_5292;
  wire CONVOLUTION_LOOP_for_for_for_asn_5294;
  wire CONVOLUTION_LOOP_for_for_for_asn_5296;
  wire CONVOLUTION_LOOP_for_for_for_asn_5298;
  wire CONVOLUTION_LOOP_for_for_for_asn_5300;
  wire CONVOLUTION_LOOP_for_for_for_asn_5302;
  wire CONVOLUTION_LOOP_for_for_for_asn_5304;
  wire CONVOLUTION_LOOP_for_for_for_asn_5306;
  wire CONVOLUTION_LOOP_for_for_for_asn_5308;
  wire CONVOLUTION_LOOP_for_for_for_asn_5310;
  wire CONVOLUTION_LOOP_for_for_for_asn_5312;
  wire CONVOLUTION_LOOP_for_for_for_asn_5314;
  wire CONVOLUTION_LOOP_for_for_for_asn_5316;
  wire CONVOLUTION_LOOP_for_for_for_asn_5318;
  wire CONVOLUTION_LOOP_for_for_for_asn_5320;
  wire CONVOLUTION_LOOP_for_for_for_asn_5322;
  wire CONVOLUTION_LOOP_for_for_for_asn_5324;
  wire CONVOLUTION_LOOP_for_for_for_asn_5326;
  wire CONVOLUTION_LOOP_for_for_for_asn_5328;
  wire CONVOLUTION_LOOP_for_for_for_asn_5330;
  wire CONVOLUTION_LOOP_for_for_for_asn_5332;
  wire CONVOLUTION_LOOP_for_for_for_asn_5334;
  wire CONVOLUTION_LOOP_for_for_for_asn_5336;
  wire CONVOLUTION_LOOP_for_for_for_asn_5338;
  wire CONVOLUTION_LOOP_for_for_for_asn_5340;
  wire CONVOLUTION_LOOP_for_for_for_asn_5342;
  wire CONVOLUTION_LOOP_for_for_for_asn_5344;
  wire CONVOLUTION_LOOP_for_for_for_asn_5346;
  wire CONVOLUTION_LOOP_for_for_for_asn_5348;
  wire CONVOLUTION_LOOP_for_for_for_asn_5350;
  wire CONVOLUTION_LOOP_for_for_for_asn_5352;
  wire CONVOLUTION_LOOP_for_for_for_asn_5354;
  wire CONVOLUTION_LOOP_for_for_for_asn_5356;
  wire CONVOLUTION_LOOP_for_for_for_asn_5358;
  wire CONVOLUTION_LOOP_for_for_for_asn_5360;
  wire CONVOLUTION_LOOP_for_for_for_asn_5362;
  wire CONVOLUTION_LOOP_for_for_for_asn_5364;
  wire CONVOLUTION_LOOP_for_for_for_asn_5366;
  wire CONVOLUTION_LOOP_for_for_for_asn_5368;
  wire CONVOLUTION_LOOP_for_for_for_asn_5370;
  wire CONVOLUTION_LOOP_for_for_for_asn_5372;
  wire CONVOLUTION_LOOP_for_for_for_asn_5374;
  wire CONVOLUTION_LOOP_for_for_for_asn_5376;
  wire CONVOLUTION_LOOP_for_for_for_asn_5378;
  wire CONVOLUTION_LOOP_for_for_for_asn_5380;
  wire CONVOLUTION_LOOP_for_for_for_asn_5382;
  wire CONVOLUTION_LOOP_for_for_for_asn_5384;
  wire CONVOLUTION_LOOP_for_for_for_asn_5386;
  wire CONVOLUTION_LOOP_for_for_for_asn_5388;
  wire CONVOLUTION_LOOP_for_for_for_asn_5390;
  wire CONVOLUTION_LOOP_for_for_for_asn_5392;
  wire CONVOLUTION_LOOP_for_for_for_asn_5394;
  wire CONVOLUTION_LOOP_for_for_for_asn_5396;
  wire CONVOLUTION_LOOP_for_for_for_asn_5398;
  wire CONVOLUTION_LOOP_for_for_for_asn_5400;
  wire CONVOLUTION_LOOP_for_for_for_asn_5402;
  wire CONVOLUTION_LOOP_for_for_for_asn_5404;
  wire CONVOLUTION_LOOP_for_for_for_asn_5406;
  wire CONVOLUTION_LOOP_for_for_for_asn_5408;
  wire CONVOLUTION_LOOP_for_for_for_asn_5410;
  wire CONVOLUTION_LOOP_for_for_for_asn_5412;
  wire CONVOLUTION_LOOP_for_for_for_asn_5414;
  wire CONVOLUTION_LOOP_for_for_for_asn_5416;
  wire CONVOLUTION_LOOP_for_for_for_asn_5418;
  wire CONVOLUTION_LOOP_for_for_for_asn_5420;
  wire CONVOLUTION_LOOP_for_for_for_asn_5422;
  wire CONVOLUTION_LOOP_for_for_for_asn_5424;
  wire CONVOLUTION_LOOP_for_for_for_asn_5426;
  wire CONVOLUTION_LOOP_for_for_for_asn_5428;
  wire CONVOLUTION_LOOP_for_for_for_asn_5430;
  wire CONVOLUTION_LOOP_for_for_for_asn_5432;
  wire CONVOLUTION_LOOP_for_for_for_asn_5434;
  wire CONVOLUTION_LOOP_for_for_for_asn_5436;
  wire CONVOLUTION_LOOP_for_for_for_asn_5438;
  wire CONVOLUTION_LOOP_for_for_for_asn_5440;
  wire CONVOLUTION_LOOP_for_for_for_asn_5442;
  wire CONVOLUTION_LOOP_for_for_for_asn_5444;
  wire CONVOLUTION_LOOP_for_for_for_asn_5446;
  wire CONVOLUTION_LOOP_for_for_for_asn_5448;
  wire CONVOLUTION_LOOP_for_for_for_asn_5450;
  wire CONVOLUTION_LOOP_for_for_for_asn_5452;
  wire CONVOLUTION_LOOP_for_for_for_asn_5454;
  wire CONVOLUTION_LOOP_for_for_for_asn_5456;
  wire CONVOLUTION_LOOP_for_for_for_asn_5458;
  wire CONVOLUTION_LOOP_for_for_for_asn_5460;
  wire CONVOLUTION_LOOP_for_for_for_asn_5462;
  wire CONVOLUTION_LOOP_for_for_for_asn_5464;
  wire CONVOLUTION_LOOP_for_for_for_asn_5466;
  wire CONVOLUTION_LOOP_for_for_for_asn_5468;
  wire CONVOLUTION_LOOP_for_for_for_asn_5470;
  wire CONVOLUTION_LOOP_for_for_for_asn_5472;
  wire CONVOLUTION_LOOP_for_for_for_asn_5474;
  wire CONVOLUTION_LOOP_for_for_for_asn_5476;
  wire CONVOLUTION_LOOP_for_for_for_asn_5478;
  wire CONVOLUTION_LOOP_for_for_for_asn_5480;
  wire CONVOLUTION_LOOP_for_for_for_asn_5482;
  wire CONVOLUTION_LOOP_for_for_for_asn_5484;
  wire CONVOLUTION_LOOP_for_for_for_asn_5486;
  wire CONVOLUTION_LOOP_for_for_for_asn_5488;
  wire CONVOLUTION_LOOP_for_for_for_asn_5490;
  wire CONVOLUTION_LOOP_for_for_for_asn_5492;
  wire CONVOLUTION_LOOP_for_for_for_asn_5494;
  wire CONVOLUTION_LOOP_for_for_for_asn_5496;
  wire CONVOLUTION_LOOP_for_for_for_asn_5498;
  wire CONVOLUTION_LOOP_for_for_for_asn_5500;
  wire CONVOLUTION_LOOP_for_for_for_asn_5502;
  wire CONVOLUTION_LOOP_for_for_for_asn_5504;
  wire CONVOLUTION_LOOP_for_for_for_asn_5506;
  wire CONVOLUTION_LOOP_for_for_for_asn_5508;
  wire CONVOLUTION_LOOP_for_for_for_asn_5510;
  wire CONVOLUTION_LOOP_for_for_for_asn_5512;
  wire and_148_rgt;
  wire PADDING_LOOP_for_row_and_1_rgt;
  wire CONVOLUTION_LOOP_for_for_for_y_and_4_rgt;
  wire CONVOLUTION_LOOP_for_for_for_y_and_2_rgt;
  wire PADDING_LOOP_chan_and_4_cse;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_10_cse;
  wire BATCH_LOOP_and_14_cse;
  reg reg_lfst_exit_STORE_LOOP_lpi_2_dfm_5_1_2_cse;
  reg reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse;
  wire PADDING_LOOP_for_for_aelse_2_and_3_cse;
  wire CONVOLUTION_LOOP_and_4_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_11_cse;
  wire and_986_cse;
  wire PADDING_LOOP_for_row_and_3_cse;
  wire CONVOLUTION_LOOP_for_for_for_for_and_12_cse;
  wire PADDING_LOOP_for_and_3_cse;
  wire PADDING_LOOP_for_for_aelse_2_and_2_cse;
  reg reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse;
  reg reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse;
  wire CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm;
  wire mux_316_itm;
  wire PADDING_LOOP_for_for_aelse_1_acc_itm_9_1;
  wire operator_8_false_2_acc_itm_4_1;
  wire operator_8_false_3_acc_itm_4_1;
  wire operator_8_false_6_acc_itm_4_1;
  wire operator_8_false_7_acc_itm_4_1;
  wire operator_8_false_8_acc_itm_3_1;
  wire operator_8_false_9_acc_itm_3_1;
  wire operator_16_false_1_acc_itm_7_1;
  wire [8:0] z_out_1_8_0;
  wire [12:0] z_out_5_12_0;
  wire [15:0] nl_z_out_5_12_0;
  wire [15:0] z_out_8_15_0;
  wire signed [24:0] nl_z_out_8_15_0;
  wire [15:0] z_out_9_15_0;
  wire signed [24:0] nl_z_out_9_15_0;
  wire [16:0] z_out_11_16_0;
  wire signed [17:0] nl_z_out_11_16_0;

  wire[0:0] mux_324_nl;
  wire[0:0] or_328_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] or_843_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl;
  wire[29:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_nl;
  wire[29:0] CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_2_nl;
  wire[31:0] PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_nl;
  wire[0:0] nor_26_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] and_788_nl;
  wire[0:0] and_789_nl;
  wire[12:0] PADDING_LOOP_for_for_index_in_acc_2_nl;
  wire[13:0] nl_PADDING_LOOP_for_for_index_in_acc_2_nl;
  wire[12:0] PADDING_LOOP_for_for_index_in_mul_2_nl;
  wire[13:0] PADDING_LOOP_for_for_index_in_mul_nl;
  wire[20:0] nl_PADDING_LOOP_for_for_index_in_mul_nl;
  wire[12:0] PADDING_LOOP_for_for_index_in_mul_1_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] and_764_nl;
  wire[0:0] nor_232_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl;
  wire[14:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl;
  wire[15:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl;
  wire[18:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl;
  wire[15:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl;
  wire[16:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl;
  wire[20:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl;
  wire[11:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_5_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] and_762_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] nor_227_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] or_603_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] and_763_nl;
  wire[0:0] nor_230_nl;
  wire[0:0] nor_187_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] or_636_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] and_790_nl;
  wire[0:0] nor_305_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] nor_296_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] nor_299_nl;
  wire[12:0] CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl;
  wire[13:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl;
  wire[12:0] CONVOLUTION_LOOP_for_for_for_index_out_mul_2_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_index_out_mul_nl;
  wire[18:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl;
  wire[15:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] nor_253_nl;
  wire[0:0] nor_255_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_249_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] and_192_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] nor_246_nl;
  wire[3:0] STORE_LOOP_mux_37_nl;
  wire[0:0] or_780_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] or_779_nl;
  wire[0:0] or_776_nl;
  wire[0:0] PADDING_LOOP_for_for_aelse_mux_nl;
  wire[0:0] BATCH_LOOP_mux_5_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] BATCH_LOOP_mux_6_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] nand_65_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] or_6_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] or_1_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] and_222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_not_2308_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] nor_389_nl;
  wire[4:0] mux_556_nl;
  wire[0:0] or_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_mux_3_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] CONVOLUTION_LOOP_mux_1_nl;
  wire[0:0] or_475_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] or_474_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_acc_and_4_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2283_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] and_917_nl;
  wire[4:0] mux_557_nl;
  wire[0:0] or_1142_nl;
  wire[0:0] PADDING_LOOP_for_for_mux_2_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] LOAD_LOOP_LOAD_LOOP_and_2_nl;
  wire[0:0] STORE_LOOP_or_2327_nl;
  wire[4:0] PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_1_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] and_915_nl;
  wire[0:0] PADDING_LOOP_PADDING_LOOP_and_2_nl;
  wire[0:0] STORE_LOOP_or_2323_nl;
  wire[0:0] and_907_nl;
  wire[0:0] and_908_nl;
  wire[0:0] and_905_nl;
  wire[0:0] and_906_nl;
  wire[0:0] STORE_LOOP_nand_nl;
  wire[0:0] STORE_LOOP_and_18_nl;
  wire[0:0] STORE_LOOP_and_25_nl;
  wire[0:0] STORE_LOOP_and_26_nl;
  wire[2:0] CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_and_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] and_913_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] STORE_LOOP_mux_31_nl;
  wire[0:0] STORE_LOOP_mux1h_2331_nl;
  wire[0:0] STORE_LOOP_mux_34_nl;
  wire[0:0] operator_42_true_1_and_nl;
  wire[0:0] STORE_LOOP_STORE_LOOP_nor_2_nl;
  wire[0:0] or_789_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2300_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2304_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2306_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2308_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2312_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2316_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2318_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2320_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2324_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2326_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2328_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2330_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2332_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2334_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2336_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2338_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2340_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2342_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2344_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2346_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2348_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2350_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2352_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2354_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2356_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2358_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2360_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2362_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2364_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2366_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2368_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2370_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2372_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2374_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2376_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2378_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2380_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2382_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2384_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2386_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2388_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2390_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2392_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2394_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2396_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2398_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2400_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2402_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2404_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2406_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2408_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2410_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2412_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2414_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2416_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2418_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2420_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2422_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2424_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2426_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2428_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2430_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2432_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2434_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2436_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2438_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2440_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2442_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2444_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2446_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2448_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2450_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2452_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2454_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2456_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2458_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2460_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2462_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2464_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2466_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2468_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2470_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2472_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2474_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2476_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2478_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2480_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2482_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2484_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2486_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2488_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2492_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2494_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2496_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2498_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2500_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2502_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2504_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2506_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2508_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2510_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2512_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2514_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2516_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2518_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2520_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2522_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2524_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2526_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2528_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2530_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2532_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2534_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2536_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2538_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2540_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2542_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2544_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2546_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2548_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2550_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2552_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2554_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2556_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2558_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2560_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2562_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2564_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2566_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2568_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2570_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2572_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2574_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2576_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2578_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2580_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2582_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2584_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2586_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2588_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2590_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2592_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2594_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2596_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2598_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2600_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2602_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2604_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2606_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2608_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2610_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2612_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2614_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2616_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2618_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2620_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2622_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2624_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2626_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2628_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2630_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2632_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2634_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2636_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2638_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2640_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2642_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2644_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2646_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2648_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2650_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2652_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2654_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2656_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2658_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2660_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2662_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2664_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2666_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2668_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2670_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2672_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2674_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2676_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2678_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2680_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2682_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2684_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2686_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2688_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2690_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2692_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2694_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2696_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2698_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2700_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2702_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2704_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2706_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2708_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2710_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2712_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2714_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2716_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2718_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2720_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2722_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2724_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2726_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2728_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2730_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2732_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2734_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2736_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2738_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2740_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2742_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2744_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2746_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2748_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2750_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2752_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2754_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2756_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2758_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2760_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2762_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2764_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2766_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2768_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2770_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2772_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2774_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2776_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2778_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2780_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2782_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2784_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2786_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2788_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2790_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2792_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2794_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2796_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2798_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2800_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2802_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2804_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2806_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2808_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2810_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2812_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2814_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2816_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2818_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2820_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2822_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2824_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2826_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2828_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2830_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2832_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2834_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2836_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2838_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2840_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2842_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2844_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2846_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2848_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2850_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2852_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2854_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2856_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2858_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2860_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2862_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2864_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2866_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2868_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2870_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2872_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2874_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2876_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2878_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2880_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2882_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2884_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2886_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2888_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2890_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2892_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2894_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2896_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2898_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2900_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2902_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2904_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2906_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2908_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2910_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2912_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2914_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2916_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2918_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2920_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2922_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2924_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2926_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2928_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2930_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2932_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2934_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2936_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2938_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2940_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2942_nl;
  wire[0:0] STORE_LOOP_mux_29_nl;
  wire[0:0] STORE_LOOP_mux_30_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl;
  wire[54:0] CONVOLUTION_LOOP_for_for_for_else_nor_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_973_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_975_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_984_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_976_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_977_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_988_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_978_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_979_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_981_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_996_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_983_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_984_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_985_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_987_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_988_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_989_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_991_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_993_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_995_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_996_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_997_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_999_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1626_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_and_nl;
  wire[9:0] PADDING_LOOP_for_for_aelse_1_acc_nl;
  wire[10:0] nl_PADDING_LOOP_for_for_aelse_1_acc_nl;
  wire[8:0] PADDING_LOOP_for_for_aelse_1_acc_1_nl;
  wire[9:0] nl_PADDING_LOOP_for_for_aelse_1_acc_1_nl;
  wire[4:0] operator_8_false_2_acc_nl;
  wire[5:0] nl_operator_8_false_2_acc_nl;
  wire[4:0] operator_8_false_3_acc_nl;
  wire[5:0] nl_operator_8_false_3_acc_nl;
  wire[0:0] PADDING_LOOP_for_mux_1_nl;
  wire[4:0] operator_8_false_6_acc_nl;
  wire[5:0] nl_operator_8_false_6_acc_nl;
  wire[4:0] operator_8_false_7_acc_nl;
  wire[5:0] nl_operator_8_false_7_acc_nl;
  wire[3:0] operator_8_false_8_acc_nl;
  wire[4:0] nl_operator_8_false_8_acc_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_not_2310_nl;
  wire[3:0] operator_8_false_9_acc_nl;
  wire[4:0] nl_operator_8_false_9_acc_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_4_nl;
  wire[0:0] CONVOLUTION_LOOP_for_mux_1_nl;
  wire[0:0] or_490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_mux_1_nl;
  wire[7:0] operator_16_false_1_acc_nl;
  wire[8:0] nl_operator_16_false_1_acc_nl;
  wire[6:0] operator_16_false_acc_nl;
  wire[7:0] nl_operator_16_false_acc_nl;
  wire[0:0] PADDING_LOOP_mux_1_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] or_639_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_and_6_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_and_7_nl;
  wire[0:0] nand_90_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] or_1104_nl;
  wire[0:0] or_334_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] or_337_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] or_376_nl;
  wire[0:0] or_375_nl;
  wire[0:0] and_130_nl;
  wire[0:0] and_129_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] or_430_nl;
  wire[0:0] or_441_nl;
  wire[0:0] or_438_nl;
  wire[0:0] nand_40_nl;
  wire[0:0] or_446_nl;
  wire[0:0] nand_43_nl;
  wire[0:0] or_524_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] nor_294_nl;
  wire[0:0] nor_295_nl;
  wire[0:0] or_546_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] or_71_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] or_70_nl;
  wire[0:0] mux_441_nl;
  wire[0:0] or_596_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] nor_272_nl;
  wire[0:0] and_165_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] nand_72_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] or_652_nl;
  wire[0:0] nand_51_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] nor_268_nl;
  wire[0:0] and_170_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] or_714_nl;
  wire[0:0] nand_54_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] or_726_nl;
  wire[0:0] or_724_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] or_380_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] nor_308_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] or_663_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] mux_506_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] or_689_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] and_139_nl;
  wire[0:0] nor_167_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] or_116_nl;
  wire[0:0] and_138_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] and_151_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] and_150_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] and_155_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] and_154_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] and_153_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] and_760_nl;
  wire[0:0] and_761_nl;
  wire[15:0] BATCH_LOOP_mux_10_nl;
  wire[15:0] BATCH_LOOP_mux_11_nl;
  wire[15:0] BATCH_LOOP_mul_3_nl;
  wire[19:0] nl_BATCH_LOOP_mul_3_nl;
  wire[15:0] dma_read_data_length_mul_5_nl;
  wire[23:0] nl_dma_read_data_length_mul_5_nl;
  wire[9:0] acc_1_nl;
  wire[10:0] nl_acc_1_nl;
  wire[8:0] operator_42_true_mux_2_nl;
  wire[7:0] operator_42_true_mux_3_nl;
  wire[0:0] operator_42_true_and_1_nl;
  wire[10:0] acc_2_nl;
  wire[11:0] nl_acc_2_nl;
  wire[8:0] else_mux_2_nl;
  wire[8:0] PADDING_LOOP_for_for_aelse_2_acc_2_nl;
  wire[9:0] nl_PADDING_LOOP_for_for_aelse_2_acc_2_nl;
  wire[0:0] else_or_1_nl;
  wire[2:0] else_else_nor_1_nl;
  wire[4:0] else_mux_3_nl;
  wire[9:0] acc_3_nl;
  wire[10:0] nl_acc_3_nl;
  wire[2:0] pad_pad_pad_nor_1_nl;
  wire[4:0] pad_mux_5_nl;
  wire[7:0] pad_mux_6_nl;
  wire[7:0] operator_8_false_mux_1_nl;
  wire[7:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_10_nl;
  wire[7:0] operator_43_true_operator_43_true_acc_1_nl;
  wire[8:0] nl_operator_43_true_operator_43_true_acc_1_nl;
  wire[0:0] operator_43_true_and_1_nl;
  wire[7:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_11_nl;
  wire[7:0] dma_read_data_length_mux_8_nl;
  wire[15:0] dma_read_data_length_mux_9_nl;
  wire[31:0] dma_read_data_length_mux_10_nl;
  wire[31:0] dma_read_data_length_mux_11_nl;
  wire[7:0] BATCH_LOOP_mux_12_nl;
  wire[15:0] BATCH_LOOP_mux_13_nl;
  wire[7:0] CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_mux1h_2_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_and_14_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_12_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_10_nl;
  wire[20:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_10_nl;
  wire[12:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_11_nl;
  wire[7:0] mux_562_nl;
  wire[7:0] dma_read_data_length_mux_12_nl;
  wire[23:0] dma_read_data_length_mux_13_nl;
  wire[23:0] LOAD_LOOP_mul_2_nl;
  wire[7:0] pad_mux_7_nl;
  wire[8:0] pad_mux_8_nl;
  wire[16:0] LOAD_LOOP_mux_2_nl;
  wire[8:0] LOAD_LOOP_mux_3_nl;
  wire[7:0] CONVOLUTION_LOOP_for_for_for_for_mux_2951_nl;
  wire[0:0] and_987_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_oswt_unreg;
  assign nl_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_oswt_unreg
      = and_dcpl_45 & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse) & (fsm_output[2]);
  wire [66:0] nl_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat;
  assign nl_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat
      = {19'b0110000000000000000 , dma_read_ctrl_rsci_idat_47_32 , 16'b0000000000000000
      , dma_read_ctrl_rsci_idat_15_0};
  wire [0:0] nl_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_oswt_unreg;
  assign nl_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_oswt_unreg
      = and_dcpl_74 & (fsm_output[2]);
  wire [66:0] nl_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat;
  assign nl_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat
      = {19'b0110000000000000000 , dma_write_ctrl_rsci_idat_47_32 , 16'b0000000000000000
      , dma_write_ctrl_rsci_idat_15_0};
  wire [0:0] nl_conv2d_cxx_catapult_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg;
  assign nl_conv2d_cxx_catapult_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg
      = and_dcpl_69 & (fsm_output[2]);
  wire [0:0] nl_conv2d_cxx_catapult_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_oswt_unreg;
  assign nl_conv2d_cxx_catapult_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_oswt_unreg
      = and_dcpl_65 & (fsm_output[2]);
  wire [63:0] nl_conv2d_cxx_catapult_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat;
  assign nl_conv2d_cxx_catapult_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat
      = {32'b11011110101011011011111011101111 , dma_write_chnl_rsci_idat_31_0};
  wire [0:0] nl_conv2d_cxx_catapult_core_plm_in_data_rsci_1_inst_plm_in_data_rsci_oswt_unreg;
  assign nl_conv2d_cxx_catapult_core_plm_in_data_rsci_1_inst_plm_in_data_rsci_oswt_unreg
      = mux_tmp_321 & and_dcpl_55 & lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1 & plm_in_data_rsci_bawt
      & lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0 & (fsm_output[2]);
  wire [0:0] nl_conv2d_cxx_catapult_core_plm_f_data_rsci_1_inst_plm_f_data_rsci_oswt_unreg;
  assign nl_conv2d_cxx_catapult_core_plm_f_data_rsci_1_inst_plm_f_data_rsci_oswt_unreg
      = mux_tmp_321 & and_dcpl_55 & lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1 & plm_f_data_rsci_bawt
      & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0) & (fsm_output[2]);
  wire [0:0] nl_conv2d_cxx_catapult_core_plm_out_data_rsci_1_inst_plm_out_data_rsci_oswt_unreg;
  assign nl_conv2d_cxx_catapult_core_plm_out_data_rsci_1_inst_plm_out_data_rsci_oswt_unreg
      = or_2_cse & and_dcpl_33 & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3 & plm_out_data_rsci_bawt
      & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0) & BATCH_LOOP_stage_v_3 & BATCH_LOOP_stage_0_4
      & (fsm_output[2]);
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_conf_info_rsci conv2d_cxx_catapult_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt(reg_conf_info_rsci_irdy_core_psct_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_ctrl_rsci conv2d_cxx_catapult_core_dma_read_ctrl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dma_read_ctrl_rsci_oswt_unreg(nl_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_oswt_unreg[0:0]),
      .dma_read_ctrl_rsci_bawt(dma_read_ctrl_rsci_bawt),
      .dma_read_ctrl_rsci_iswt0(reg_dma_read_ctrl_rsci_ivld_core_psct_cse),
      .dma_read_ctrl_rsci_irdy_mxwt(dma_read_ctrl_rsci_irdy_mxwt),
      .dma_read_ctrl_rsci_idat(nl_conv2d_cxx_catapult_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat[66:0])
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_ctrl_rsci conv2d_cxx_catapult_core_dma_write_ctrl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .core_wen(core_wen),
      .dma_write_ctrl_rsci_oswt_unreg(nl_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_oswt_unreg[0:0]),
      .dma_write_ctrl_rsci_bawt(dma_write_ctrl_rsci_bawt),
      .dma_write_ctrl_rsci_iswt0(reg_dma_write_ctrl_rsci_ivld_core_psct_cse),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_ctrl_rsci_idat(nl_conv2d_cxx_catapult_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat[66:0])
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_read_chnl_rsci conv2d_cxx_catapult_core_dma_read_chnl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .core_wen(core_wen),
      .dma_read_chnl_rsci_oswt_unreg(nl_conv2d_cxx_catapult_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg[0:0]),
      .dma_read_chnl_rsci_bawt(dma_read_chnl_rsci_bawt),
      .dma_read_chnl_rsci_iswt0(reg_dma_read_chnl_rsci_irdy_core_psct_cse),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .dma_read_chnl_rsci_idat_mxwt(dma_read_chnl_rsci_idat_mxwt)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_dma_write_chnl_rsci conv2d_cxx_catapult_core_dma_write_chnl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .core_wen(core_wen),
      .dma_write_chnl_rsci_oswt_unreg(nl_conv2d_cxx_catapult_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_oswt_unreg[0:0]),
      .dma_write_chnl_rsci_bawt(dma_write_chnl_rsci_bawt),
      .dma_write_chnl_rsci_iswt0(reg_dma_write_chnl_rsci_ivld_core_psct_cse),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .dma_write_chnl_rsci_idat(nl_conv2d_cxx_catapult_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat[63:0])
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_acc_done_rsci conv2d_cxx_catapult_core_acc_done_rsci_inst
      (
      .acc_done_rsc_vld(acc_done_rsc_vld),
      .core_wten(core_wten),
      .acc_done_rsci_iswt0(reg_acc_done_rsci_ivld_core_psct_cse)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_in_data_rsci_1 conv2d_cxx_catapult_core_plm_in_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_data_rsci_q_d(plm_in_data_rsci_q_d),
      .plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_in_data_rsci_oswt_unreg(nl_conv2d_cxx_catapult_core_plm_in_data_rsci_1_inst_plm_in_data_rsci_oswt_unreg[0:0]),
      .plm_in_data_rsci_bawt(plm_in_data_rsci_bawt),
      .plm_in_data_rsci_iswt0(reg_plm_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse),
      .plm_in_data_rsci_oswt_unreg_1(and_257_rmff),
      .plm_in_data_rsci_iswt0_1(reg_plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .plm_in_data_rsci_q_d_mxwt(plm_in_data_rsci_q_d_mxwt),
      .plm_in_data_rsci_we_d_pff(plm_in_data_rsci_we_d_iff),
      .plm_in_data_rsci_iswt0_pff(and_261_rmff),
      .plm_in_data_rsci_iswt0_1_pff(and_253_rmff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_f_data_rsci_1 conv2d_cxx_catapult_core_plm_f_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_f_data_rsci_q_d(plm_f_data_rsci_q_d),
      .plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_f_data_rsci_oswt_unreg(nl_conv2d_cxx_catapult_core_plm_f_data_rsci_1_inst_plm_f_data_rsci_oswt_unreg[0:0]),
      .plm_f_data_rsci_bawt(plm_f_data_rsci_bawt),
      .plm_f_data_rsci_iswt0(reg_plm_f_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse),
      .plm_f_data_rsci_oswt_unreg_1(and_257_rmff),
      .plm_f_data_rsci_iswt0_1(reg_plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .plm_f_data_rsci_q_d_mxwt(plm_f_data_rsci_q_d_mxwt),
      .plm_f_data_rsci_we_d_pff(plm_f_data_rsci_we_d_iff),
      .plm_f_data_rsci_iswt0_pff(and_255_rmff),
      .plm_f_data_rsci_iswt0_1_pff(and_253_rmff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_plm_out_data_rsci_1 conv2d_cxx_catapult_core_plm_out_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_data_rsci_q_d(plm_out_data_rsci_q_d),
      .plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_out_data_rsci_oswt_unreg(nl_conv2d_cxx_catapult_core_plm_out_data_rsci_1_inst_plm_out_data_rsci_oswt_unreg[0:0]),
      .plm_out_data_rsci_bawt(plm_out_data_rsci_bawt),
      .plm_out_data_rsci_iswt0(reg_plm_out_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse),
      .plm_out_data_rsci_oswt_unreg_1(or_tmp_676),
      .plm_out_data_rsci_iswt0_1(reg_plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .plm_out_data_rsci_q_d_mxwt(plm_out_data_rsci_q_d_mxwt),
      .plm_out_data_rsci_we_d_pff(plm_out_data_rsci_we_d_iff),
      .plm_out_data_rsci_iswt0_pff(and_247_rmff),
      .plm_out_data_rsci_iswt0_1_pff(and_245_rmff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_staller conv2d_cxx_catapult_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_fsm conv2d_cxx_catapult_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output),
      .BATCH_LOOP_C_0_tr0(and_dcpl_16)
    );
  assign or_328_nl = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (operator_8_false_4_acc_tmp[8:3]!=6'b000000)
      | mux_376_cse;
  assign mux_324_nl = MUX_s_1_2_2(mux_376_cse, or_328_nl, operator_8_false_9_acc_itm_3_1);
  assign nand_25_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_240_cse
      | (operator_8_false_4_acc_tmp[8:3]!=6'b000000) | mux_376_cse)));
  assign mux_325_cse = MUX_s_1_2_2(mux_324_nl, nand_25_nl, operator_8_false_8_acc_itm_3_1);
  assign nor_291_cse = ~(and_769_cse | and_770_cse | mux_325_cse);
  assign BATCH_LOOP_and_cse = core_wen & (fsm_output[2]) & or_316_cse & or_453_cse
      & nor_291_cse & BATCH_LOOP_and_6_tmp;
  assign LOAD_CTRL_LOOP_and_cse = core_wen & (fsm_output[2]) & mux_tmp_319 & BATCH_LOOP_and_6_tmp;
  assign and_245_rmff = mux_tmp_321 & and_dcpl_23 & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1)
      & lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0 & (fsm_output[2]);
  assign and_247_rmff = mux_tmp_321 & and_dcpl_22 & lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2
      & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1) & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0)
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_2 & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2
      & (fsm_output[2]);
  assign and_253_rmff = and_dcpl_45 & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse
      & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse) & (fsm_output[2]);
  assign and_255_rmff = and_dcpl_48 & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse)
      & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse) & (fsm_output[2]);
  assign and_257_rmff = mux_tmp_321 & and_dcpl_23 & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1)
      & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0) & (fsm_output[2]);
  assign and_261_rmff = and_dcpl_48 & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse)
      & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse & (fsm_output[2]);
  assign CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff = MUX_v_14_2_2(CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2,
      plm_out_data_rsci_wadr_d_reg, or_tmp_709);
  assign or_843_nl = (~ (fsm_output[2])) | (~ mux_tmp_321) | not_tmp_164 | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2)
      | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1 | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0);
  assign CONVOLUTION_LOOP_for_for_for_index_out_mux_1_rmff = MUX_v_14_2_2(CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2,
      plm_out_data_rsci_radr_d_reg, or_843_nl);
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl = MUX_s_1_324_2(buf_acc_data_0_0_0_sva_dfm_mx0,
      buf_acc_data_0_1_0_sva_dfm_mx0, buf_acc_data_0_2_0_sva_dfm_mx0, buf_acc_data_0_3_0_sva_dfm_mx0,
      buf_acc_data_0_4_0_sva_dfm_mx0, buf_acc_data_0_5_0_sva_dfm_mx0, buf_acc_data_0_6_0_sva_dfm_mx0,
      buf_acc_data_0_7_0_sva_dfm_mx0, buf_acc_data_0_8_0_sva_dfm_mx0, buf_acc_data_0_9_0_sva_dfm_mx0,
      buf_acc_data_0_10_0_sva_dfm_mx0, buf_acc_data_0_11_0_sva_dfm_mx0, buf_acc_data_0_12_0_sva_dfm_mx0,
      buf_acc_data_0_13_0_sva_dfm_mx0, buf_acc_data_0_14_0_sva_dfm_mx0, buf_acc_data_0_15_0_sva_dfm_mx0,
      buf_acc_data_0_16_0_sva_dfm_mx0, buf_acc_data_0_17_0_sva_dfm_mx0, buf_acc_data_1_0_0_sva_dfm_mx0,
      buf_acc_data_1_1_0_sva_dfm_mx0, buf_acc_data_1_2_0_sva_dfm_mx0, buf_acc_data_1_3_0_sva_dfm_mx0,
      buf_acc_data_1_4_0_sva_dfm_mx0, buf_acc_data_1_5_0_sva_dfm_mx0, buf_acc_data_1_6_0_sva_dfm_mx0,
      buf_acc_data_1_7_0_sva_dfm_mx0, buf_acc_data_1_8_0_sva_dfm_mx0, buf_acc_data_1_9_0_sva_dfm_mx0,
      buf_acc_data_1_10_0_sva_dfm_mx0, buf_acc_data_1_11_0_sva_dfm_mx0, buf_acc_data_1_12_0_sva_dfm_mx0,
      buf_acc_data_1_13_0_sva_dfm_mx0, buf_acc_data_1_14_0_sva_dfm_mx0, buf_acc_data_1_15_0_sva_dfm_mx0,
      buf_acc_data_1_16_0_sva_dfm_mx0, buf_acc_data_1_17_0_sva_dfm_mx0, buf_acc_data_2_0_0_sva_dfm_mx0,
      buf_acc_data_2_1_0_sva_dfm_mx0, buf_acc_data_2_2_0_sva_dfm_mx0, buf_acc_data_2_3_0_sva_dfm_mx0,
      buf_acc_data_2_4_0_sva_dfm_mx0, buf_acc_data_2_5_0_sva_dfm_mx0, buf_acc_data_2_6_0_sva_dfm_mx0,
      buf_acc_data_2_7_0_sva_dfm_mx0, buf_acc_data_2_8_0_sva_dfm_mx0, buf_acc_data_2_9_0_sva_dfm_mx0,
      buf_acc_data_2_10_0_sva_dfm_mx0, buf_acc_data_2_11_0_sva_dfm_mx0, buf_acc_data_2_12_0_sva_dfm_mx0,
      buf_acc_data_2_13_0_sva_dfm_mx0, buf_acc_data_2_14_0_sva_dfm_mx0, buf_acc_data_2_15_0_sva_dfm_mx0,
      buf_acc_data_2_16_0_sva_dfm_mx0, buf_acc_data_2_17_0_sva_dfm_mx0, buf_acc_data_3_0_0_sva_dfm_mx0,
      buf_acc_data_3_1_0_sva_dfm_mx0, buf_acc_data_3_2_0_sva_dfm_mx0, buf_acc_data_3_3_0_sva_dfm_mx0,
      buf_acc_data_3_4_0_sva_dfm_mx0, buf_acc_data_3_5_0_sva_dfm_mx0, buf_acc_data_3_6_0_sva_dfm_mx0,
      buf_acc_data_3_7_0_sva_dfm_mx0, buf_acc_data_3_8_0_sva_dfm_mx0, buf_acc_data_3_9_0_sva_dfm_mx0,
      buf_acc_data_3_10_0_sva_dfm_mx0, buf_acc_data_3_11_0_sva_dfm_mx0, buf_acc_data_3_12_0_sva_dfm_mx0,
      buf_acc_data_3_13_0_sva_dfm_mx0, buf_acc_data_3_14_0_sva_dfm_mx0, buf_acc_data_3_15_0_sva_dfm_mx0,
      buf_acc_data_3_16_0_sva_dfm_mx0, buf_acc_data_3_17_0_sva_dfm_mx0, buf_acc_data_4_0_0_sva_dfm_mx0,
      buf_acc_data_4_1_0_sva_dfm_mx0, buf_acc_data_4_2_0_sva_dfm_mx0, buf_acc_data_4_3_0_sva_dfm_mx0,
      buf_acc_data_4_4_0_sva_dfm_mx0, buf_acc_data_4_5_0_sva_dfm_mx0, buf_acc_data_4_6_0_sva_dfm_mx0,
      buf_acc_data_4_7_0_sva_dfm_mx0, buf_acc_data_4_8_0_sva_dfm_mx0, buf_acc_data_4_9_0_sva_dfm_mx0,
      buf_acc_data_4_10_0_sva_dfm_mx0, buf_acc_data_4_11_0_sva_dfm_mx0, buf_acc_data_4_12_0_sva_dfm_mx0,
      buf_acc_data_4_13_0_sva_dfm_mx0, buf_acc_data_4_14_0_sva_dfm_mx0, buf_acc_data_4_15_0_sva_dfm_mx0,
      buf_acc_data_4_16_0_sva_dfm_mx0, buf_acc_data_4_17_0_sva_dfm_mx0, buf_acc_data_5_0_0_sva_dfm_mx0,
      buf_acc_data_5_1_0_sva_dfm_mx0, buf_acc_data_5_2_0_sva_dfm_mx0, buf_acc_data_5_3_0_sva_dfm_mx0,
      buf_acc_data_5_4_0_sva_dfm_mx0, buf_acc_data_5_5_0_sva_dfm_mx0, buf_acc_data_5_6_0_sva_dfm_mx0,
      buf_acc_data_5_7_0_sva_dfm_mx0, buf_acc_data_5_8_0_sva_dfm_mx0, buf_acc_data_5_9_0_sva_dfm_mx0,
      buf_acc_data_5_10_0_sva_dfm_mx0, buf_acc_data_5_11_0_sva_dfm_mx0, buf_acc_data_5_12_0_sva_dfm_mx0,
      buf_acc_data_5_13_0_sva_dfm_mx0, buf_acc_data_5_14_0_sva_dfm_mx0, buf_acc_data_5_15_0_sva_dfm_mx0,
      buf_acc_data_5_16_0_sva_dfm_mx0, buf_acc_data_5_17_0_sva_dfm_mx0, buf_acc_data_6_0_0_sva_dfm_mx0,
      buf_acc_data_6_1_0_sva_dfm_mx0, buf_acc_data_6_2_0_sva_dfm_mx0, buf_acc_data_6_3_0_sva_dfm_mx0,
      buf_acc_data_6_4_0_sva_dfm_mx0, buf_acc_data_6_5_0_sva_dfm_mx0, buf_acc_data_6_6_0_sva_dfm_mx0,
      buf_acc_data_6_7_0_sva_dfm_mx0, buf_acc_data_6_8_0_sva_dfm_mx0, buf_acc_data_6_9_0_sva_dfm_mx0,
      buf_acc_data_6_10_0_sva_dfm_mx0, buf_acc_data_6_11_0_sva_dfm_mx0, buf_acc_data_6_12_0_sva_dfm_mx0,
      buf_acc_data_6_13_0_sva_dfm_mx0, buf_acc_data_6_14_0_sva_dfm_mx0, buf_acc_data_6_15_0_sva_dfm_mx0,
      buf_acc_data_6_16_0_sva_dfm_mx0, buf_acc_data_6_17_0_sva_dfm_mx0, buf_acc_data_7_0_0_sva_dfm_mx0,
      buf_acc_data_7_1_0_sva_dfm_mx0, buf_acc_data_7_2_0_sva_dfm_mx0, buf_acc_data_7_3_0_sva_dfm_mx0,
      buf_acc_data_7_4_0_sva_dfm_mx0, buf_acc_data_7_5_0_sva_dfm_mx0, buf_acc_data_7_6_0_sva_dfm_mx0,
      buf_acc_data_7_7_0_sva_dfm_mx0, buf_acc_data_7_8_0_sva_dfm_mx0, buf_acc_data_7_9_0_sva_dfm_mx0,
      buf_acc_data_7_10_0_sva_dfm_mx0, buf_acc_data_7_11_0_sva_dfm_mx0, buf_acc_data_7_12_0_sva_dfm_mx0,
      buf_acc_data_7_13_0_sva_dfm_mx0, buf_acc_data_7_14_0_sva_dfm_mx0, buf_acc_data_7_15_0_sva_dfm_mx0,
      buf_acc_data_7_16_0_sva_dfm_mx0, buf_acc_data_7_17_0_sva_dfm_mx0, buf_acc_data_8_0_0_sva_dfm_mx0,
      buf_acc_data_8_1_0_sva_dfm_mx0, buf_acc_data_8_2_0_sva_dfm_mx0, buf_acc_data_8_3_0_sva_dfm_mx0,
      buf_acc_data_8_4_0_sva_dfm_mx0, buf_acc_data_8_5_0_sva_dfm_mx0, buf_acc_data_8_6_0_sva_dfm_mx0,
      buf_acc_data_8_7_0_sva_dfm_mx0, buf_acc_data_8_8_0_sva_dfm_mx0, buf_acc_data_8_9_0_sva_dfm_mx0,
      buf_acc_data_8_10_0_sva_dfm_mx0, buf_acc_data_8_11_0_sva_dfm_mx0, buf_acc_data_8_12_0_sva_dfm_mx0,
      buf_acc_data_8_13_0_sva_dfm_mx0, buf_acc_data_8_14_0_sva_dfm_mx0, buf_acc_data_8_15_0_sva_dfm_mx0,
      buf_acc_data_8_16_0_sva_dfm_mx0, buf_acc_data_8_17_0_sva_dfm_mx0, buf_acc_data_9_0_0_sva_dfm_mx0,
      buf_acc_data_9_1_0_sva_dfm_mx0, buf_acc_data_9_2_0_sva_dfm_mx0, buf_acc_data_9_3_0_sva_dfm_mx0,
      buf_acc_data_9_4_0_sva_dfm_mx0, buf_acc_data_9_5_0_sva_dfm_mx0, buf_acc_data_9_6_0_sva_dfm_mx0,
      buf_acc_data_9_7_0_sva_dfm_mx0, buf_acc_data_9_8_0_sva_dfm_mx0, buf_acc_data_9_9_0_sva_dfm_mx0,
      buf_acc_data_9_10_0_sva_dfm_mx0, buf_acc_data_9_11_0_sva_dfm_mx0, buf_acc_data_9_12_0_sva_dfm_mx0,
      buf_acc_data_9_13_0_sva_dfm_mx0, buf_acc_data_9_14_0_sva_dfm_mx0, buf_acc_data_9_15_0_sva_dfm_mx0,
      buf_acc_data_9_16_0_sva_dfm_mx0, buf_acc_data_9_17_0_sva_dfm_mx0, buf_acc_data_10_0_0_sva_dfm_mx0,
      buf_acc_data_10_1_0_sva_dfm_mx0, buf_acc_data_10_2_0_sva_dfm_mx0, buf_acc_data_10_3_0_sva_dfm_mx0,
      buf_acc_data_10_4_0_sva_dfm_mx0, buf_acc_data_10_5_0_sva_dfm_mx0, buf_acc_data_10_6_0_sva_dfm_mx0,
      buf_acc_data_10_7_0_sva_dfm_mx0, buf_acc_data_10_8_0_sva_dfm_mx0, buf_acc_data_10_9_0_sva_dfm_mx0,
      buf_acc_data_10_10_0_sva_dfm_mx0, buf_acc_data_10_11_0_sva_dfm_mx0, buf_acc_data_10_12_0_sva_dfm_mx0,
      buf_acc_data_10_13_0_sva_dfm_mx0, buf_acc_data_10_14_0_sva_dfm_mx0, buf_acc_data_10_15_0_sva_dfm_mx0,
      buf_acc_data_10_16_0_sva_dfm_mx0, buf_acc_data_10_17_0_sva_dfm_mx0, buf_acc_data_11_0_0_sva_dfm_mx0,
      buf_acc_data_11_1_0_sva_dfm_mx0, buf_acc_data_11_2_0_sva_dfm_mx0, buf_acc_data_11_3_0_sva_dfm_mx0,
      buf_acc_data_11_4_0_sva_dfm_mx0, buf_acc_data_11_5_0_sva_dfm_mx0, buf_acc_data_11_6_0_sva_dfm_mx0,
      buf_acc_data_11_7_0_sva_dfm_mx0, buf_acc_data_11_8_0_sva_dfm_mx0, buf_acc_data_11_9_0_sva_dfm_mx0,
      buf_acc_data_11_10_0_sva_dfm_mx0, buf_acc_data_11_11_0_sva_dfm_mx0, buf_acc_data_11_12_0_sva_dfm_mx0,
      buf_acc_data_11_13_0_sva_dfm_mx0, buf_acc_data_11_14_0_sva_dfm_mx0, buf_acc_data_11_15_0_sva_dfm_mx0,
      buf_acc_data_11_16_0_sva_dfm_mx0, buf_acc_data_11_17_0_sva_dfm_mx0, buf_acc_data_12_0_0_sva_dfm_mx0,
      buf_acc_data_12_1_0_sva_dfm_mx0, buf_acc_data_12_2_0_sva_dfm_mx0, buf_acc_data_12_3_0_sva_dfm_mx0,
      buf_acc_data_12_4_0_sva_dfm_mx0, buf_acc_data_12_5_0_sva_dfm_mx0, buf_acc_data_12_6_0_sva_dfm_mx0,
      buf_acc_data_12_7_0_sva_dfm_mx0, buf_acc_data_12_8_0_sva_dfm_mx0, buf_acc_data_12_9_0_sva_dfm_mx0,
      buf_acc_data_12_10_0_sva_dfm_mx0, buf_acc_data_12_11_0_sva_dfm_mx0, buf_acc_data_12_12_0_sva_dfm_mx0,
      buf_acc_data_12_13_0_sva_dfm_mx0, buf_acc_data_12_14_0_sva_dfm_mx0, buf_acc_data_12_15_0_sva_dfm_mx0,
      buf_acc_data_12_16_0_sva_dfm_mx0, buf_acc_data_12_17_0_sva_dfm_mx0, buf_acc_data_13_0_0_sva_dfm_mx0,
      buf_acc_data_13_1_0_sva_dfm_mx0, buf_acc_data_13_2_0_sva_dfm_mx0, buf_acc_data_13_3_0_sva_dfm_mx0,
      buf_acc_data_13_4_0_sva_dfm_mx0, buf_acc_data_13_5_0_sva_dfm_mx0, buf_acc_data_13_6_0_sva_dfm_mx0,
      buf_acc_data_13_7_0_sva_dfm_mx0, buf_acc_data_13_8_0_sva_dfm_mx0, buf_acc_data_13_9_0_sva_dfm_mx0,
      buf_acc_data_13_10_0_sva_dfm_mx0, buf_acc_data_13_11_0_sva_dfm_mx0, buf_acc_data_13_12_0_sva_dfm_mx0,
      buf_acc_data_13_13_0_sva_dfm_mx0, buf_acc_data_13_14_0_sva_dfm_mx0, buf_acc_data_13_15_0_sva_dfm_mx0,
      buf_acc_data_13_16_0_sva_dfm_mx0, buf_acc_data_13_17_0_sva_dfm_mx0, buf_acc_data_14_0_0_sva_dfm_mx0,
      buf_acc_data_14_1_0_sva_dfm_mx0, buf_acc_data_14_2_0_sva_dfm_mx0, buf_acc_data_14_3_0_sva_dfm_mx0,
      buf_acc_data_14_4_0_sva_dfm_mx0, buf_acc_data_14_5_0_sva_dfm_mx0, buf_acc_data_14_6_0_sva_dfm_mx0,
      buf_acc_data_14_7_0_sva_dfm_mx0, buf_acc_data_14_8_0_sva_dfm_mx0, buf_acc_data_14_9_0_sva_dfm_mx0,
      buf_acc_data_14_10_0_sva_dfm_mx0, buf_acc_data_14_11_0_sva_dfm_mx0, buf_acc_data_14_12_0_sva_dfm_mx0,
      buf_acc_data_14_13_0_sva_dfm_mx0, buf_acc_data_14_14_0_sva_dfm_mx0, buf_acc_data_14_15_0_sva_dfm_mx0,
      buf_acc_data_14_16_0_sva_dfm_mx0, buf_acc_data_14_17_0_sva_dfm_mx0, buf_acc_data_15_0_0_sva_dfm_mx0,
      buf_acc_data_15_1_0_sva_dfm_mx0, buf_acc_data_15_2_0_sva_dfm_mx0, buf_acc_data_15_3_0_sva_dfm_mx0,
      buf_acc_data_15_4_0_sva_dfm_mx0, buf_acc_data_15_5_0_sva_dfm_mx0, buf_acc_data_15_6_0_sva_dfm_mx0,
      buf_acc_data_15_7_0_sva_dfm_mx0, buf_acc_data_15_8_0_sva_dfm_mx0, buf_acc_data_15_9_0_sva_dfm_mx0,
      buf_acc_data_15_10_0_sva_dfm_mx0, buf_acc_data_15_11_0_sva_dfm_mx0, buf_acc_data_15_12_0_sva_dfm_mx0,
      buf_acc_data_15_13_0_sva_dfm_mx0, buf_acc_data_15_14_0_sva_dfm_mx0, buf_acc_data_15_15_0_sva_dfm_mx0,
      buf_acc_data_15_16_0_sva_dfm_mx0, buf_acc_data_15_17_0_sva_dfm_mx0, buf_acc_data_16_0_0_sva_dfm_mx0,
      buf_acc_data_16_1_0_sva_dfm_mx0, buf_acc_data_16_2_0_sva_dfm_mx0, buf_acc_data_16_3_0_sva_dfm_mx0,
      buf_acc_data_16_4_0_sva_dfm_mx0, buf_acc_data_16_5_0_sva_dfm_mx0, buf_acc_data_16_6_0_sva_dfm_mx0,
      buf_acc_data_16_7_0_sva_dfm_mx0, buf_acc_data_16_8_0_sva_dfm_mx0, buf_acc_data_16_9_0_sva_dfm_mx0,
      buf_acc_data_16_10_0_sva_dfm_mx0, buf_acc_data_16_11_0_sva_dfm_mx0, buf_acc_data_16_12_0_sva_dfm_mx0,
      buf_acc_data_16_13_0_sva_dfm_mx0, buf_acc_data_16_14_0_sva_dfm_mx0, buf_acc_data_16_15_0_sva_dfm_mx0,
      buf_acc_data_16_16_0_sva_dfm_mx0, buf_acc_data_16_17_0_sva_dfm_mx0, buf_acc_data_17_0_0_sva_dfm_mx0,
      buf_acc_data_17_1_0_sva_dfm_mx0, buf_acc_data_17_2_0_sva_dfm_mx0, buf_acc_data_17_3_0_sva_dfm_mx0,
      buf_acc_data_17_4_0_sva_dfm_mx0, buf_acc_data_17_5_0_sva_dfm_mx0, buf_acc_data_17_6_0_sva_dfm_mx0,
      buf_acc_data_17_7_0_sva_dfm_mx0, buf_acc_data_17_8_0_sva_dfm_mx0, buf_acc_data_17_9_0_sva_dfm_mx0,
      buf_acc_data_17_10_0_sva_dfm_mx0, buf_acc_data_17_11_0_sva_dfm_mx0, buf_acc_data_17_12_0_sva_dfm_mx0,
      buf_acc_data_17_13_0_sva_dfm_mx0, buf_acc_data_17_14_0_sva_dfm_mx0, buf_acc_data_17_15_0_sva_dfm_mx0,
      buf_acc_data_17_16_0_sva_dfm_mx0, buf_acc_data_17_17_0_sva_dfm_mx0, {CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_2
      , CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_2
      , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0});
  assign CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_1_nl
      = ~((~(CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl | CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1))
      | CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_1_nl,
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5,
      or_tmp_709);
  assign CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl = ~(MUX_v_30_2_2((CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_45_1_1[29:0]),
      30'b111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_nl
      = ~(MUX_v_30_2_2(CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl, 30'b111111111111111111111111111111,
      CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff = MUX_v_30_2_2(CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_nl,
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4,
      or_tmp_709);
  assign CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_2_nl
      = ~((~((CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_45_1_1[30])
      | CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_5_rmff = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_2_nl,
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3,
      or_tmp_709);
  assign LOAD_LOOP_i_mux_rmff = MUX_v_16_2_2(LOAD_LOOP_i_lpi_2, plm_f_data_rsci_wadr_d_reg,
      or_tmp_714);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff = MUX_v_16_2_2(CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1,
      plm_f_data_rsci_radr_d_reg, or_tmp_715);
  assign LOAD_LOOP_data_ac_mux_rmff = MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
      plm_f_data_rsci_d_d_reg, or_tmp_714);
  assign PADDING_LOOP_for_for_index_in_mux_rmff = MUX_v_14_2_2(PADDING_LOOP_for_for_index_in_acc_itm_1,
      plm_in_data_rsci_wadr_d_reg, or_tmp_717);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff = MUX_v_14_2_2(CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1,
      plm_in_data_rsci_radr_d_reg, or_tmp_715);
  assign PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      dma_read_chnl_rsci_idat_mxwt, PADDING_LOOP_for_for_land_2_lpi_2_dfm_1);
  assign PADDING_LOOP_for_for_mux_rmff = MUX_v_32_2_2(PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_nl,
      plm_in_data_rsci_d_d_reg, or_tmp_717);
  assign STORE_LOOP_and_703_cse = core_wen & (fsm_output[2]) & BATCH_LOOP_and_4_tmp;
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_cse = core_wen & (~((~ (fsm_output[2]))
      | or_dcpl_56));
  assign STORE_LOOP_and_709_cse = core_wen & (~((~ (fsm_output[2])) | (~ mux_tmp_352)
      | nand_109_cse));
  assign and_830_cse = exit_BATCH_LOOP_lpi_2_dfm_2_1 & exitL_exit_STORE_LOOP_sva;
  assign or_81_cse = lfst_exit_STORE_LOOP_lpi_2_1 | (~ lfst_exit_STORE_LOOP_lpi_2_0)
      | (~ lfst_exit_STORE_LOOP_lpi_2_2) | exitL_exit_STORE_LOOP_sva;
  assign PADDING_LOOP_chan_and_cse = core_wen & ((fsm_output[3:2]!=2'b00));
  assign PADDING_LOOP_chan_and_4_cse = PADDING_LOOP_chan_and_cse & ((~ or_dcpl_60)
      | (fsm_output[3]));
  assign or_1066_cse = (~ CONVOLUTION_LOOP_for_for_if_equal_tmp) | (operator_8_false_8_acc_tmp[8:5]!=4'b0000);
  assign and_769_cse = or_1066_cse & operator_8_false_6_acc_itm_4_1;
  assign or_1067_cse = (~ CONVOLUTION_LOOP_for_for_for_if_2_equal_tmp) | (operator_8_false_7_acc_tmp[8:5]!=4'b0000);
  assign and_770_cse = or_1067_cse & operator_8_false_7_acc_itm_4_1;
  assign nor_240_cse = ~((~ operator_8_false_9_acc_itm_3_1) | CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp);
  assign or_453_cse = (~((~ CONVOLUTION_LOOP_for_for_for_if_1_equal_cse) | (z_out_4[8:5]!=4'b0000)))
      | (CONVOLUTION_LOOP_for_acc_tmp[5]);
  assign or_324_cse = or_tmp_293 | and_830_cse;
  assign nor_26_nl = ~(BATCH_LOOP_asn_itm_1 | (~ BATCH_LOOP_and_4_tmp));
  assign mux_376_cse = MUX_s_1_2_2(or_156_cse, or_324_cse, nor_26_nl);
  assign or_1062_cse = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (operator_8_false_4_acc_tmp[8:3]!=6'b000000);
  assign and_765_cse = or_1062_cse & operator_8_false_9_acc_itm_3_1;
  assign and_788_nl = STORE_LOOP_or_2335_tmp & or_tmp_440;
  assign and_789_nl = lfst_exit_STORE_LOOP_lpi_2_1 & or_tmp_440;
  assign mux_377_nl = MUX_s_1_2_2(and_788_nl, and_789_nl, or_214_cse);
  assign PADDING_LOOP_for_for_aelse_2_and_2_cse = core_wen & mux_377_nl & BATCH_LOOP_and_6_tmp
      & (fsm_output[2]);
  assign or_214_cse = (~ BATCH_LOOP_and_4_tmp) | BATCH_LOOP_asn_itm_1;
  assign nor_93_cse = ~(STORE_LOOP_or_2335_tmp | (~ STORE_LOOP_STORE_LOOP_or_tmp));
  assign nor_90_cse = ~(lfst_exit_STORE_LOOP_lpi_2_1 | (~ lfst_exit_STORE_LOOP_lpi_2_2));
  assign and_148_rgt = or_214_cse & (~ lfst_exit_STORE_LOOP_lpi_2_0) & BATCH_LOOP_and_6_tmp
      & (fsm_output[2]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_10_cse = core_wen & (~ or_dcpl_73)
      & (fsm_output[2]);
  assign mux_430_nl = MUX_s_1_2_2(mux_tmp_421, or_tmp_492, and_830_cse);
  assign nor_27_nl = ~(STORE_LOOP_or_2335_tmp | (~ STORE_LOOP_or_2336_tmp) | (~ STORE_LOOP_STORE_LOOP_or_tmp));
  assign mux_431_nl = MUX_s_1_2_2(or_tmp_492, mux_430_nl, nor_27_nl);
  assign mux_429_nl = MUX_s_1_2_2(mux_tmp_421, or_tmp_492, or_81_cse);
  assign mux_432_nl = MUX_s_1_2_2(mux_431_nl, mux_429_nl, or_214_cse);
  assign BATCH_LOOP_and_14_cse = core_wen & mux_432_nl & BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign BATCH_LOOP_and_10_cse = core_wen & (fsm_output[2]) & BATCH_LOOP_and_6_tmp;
  assign STORE_LOOP_and_30_cse = exit_LOAD_LOOP_lpi_2_dfm_1 & STORE_LOOP_equal_tmp_6;
  assign STORE_LOOP_and_32_cse = exit_PADDING_LOOP_lpi_2_dfm_3 & STORE_LOOP_equal_tmp_5;
  assign STORE_LOOP_and_33_cse = (~ exit_CONVOLUTION_LOOP_lpi_2_dfm_2_mx0w0) & STORE_LOOP_equal_tmp_2_mx0w0;
  assign STORE_LOOP_and_29_cse = (~ exit_LOAD_LOOP_lpi_2_dfm_1) & STORE_LOOP_equal_tmp_6;
  assign STORE_LOOP_and_31_cse = (~ exit_PADDING_LOOP_lpi_2_dfm_3) & STORE_LOOP_equal_tmp_5;
  assign nor_229_cse = ~((~ operator_8_false_8_acc_itm_3_1) | CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp);
  assign PADDING_LOOP_for_for_aelse_2_and_1_cse = core_wen & (fsm_output[2]);
  assign PADDING_LOOP_for_for_aelse_2_and_3_cse = PADDING_LOOP_for_for_aelse_2_and_1_cse
      & (~(mux_tmp_356 | (~ BATCH_LOOP_and_6_tmp)));
  assign CONVOLUTION_LOOP_and_4_cse = PADDING_LOOP_for_for_aelse_2_and_1_cse & (~
      or_dcpl_85);
  assign and_790_nl = (~(nor_303_cse | STORE_LOOP_or_2335_tmp | STORE_LOOP_or_2336_tmp
      | (~ STORE_LOOP_STORE_LOOP_or_tmp))) & (~(and_830_cse | mux_tmp_472));
  assign nor_305_nl = ~(nor_306_cse | lfst_exit_STORE_LOOP_lpi_2_1 | lfst_exit_STORE_LOOP_lpi_2_0
      | (~ lfst_exit_STORE_LOOP_lpi_2_2) | exitL_exit_STORE_LOOP_sva | mux_tmp_472);
  assign mux_480_nl = MUX_s_1_2_2(and_790_nl, nor_305_nl, or_214_cse);
  assign CONVOLUTION_LOOP_for_for_for_else_and_836_cse = core_wen & ((mux_480_nl
      & BATCH_LOOP_and_6_tmp & (fsm_output[2])) | or_tmp_801);
  assign nor_300_nl = ~(STORE_LOOP_or_2335_tmp | STORE_LOOP_or_2336_tmp | (~ STORE_LOOP_STORE_LOOP_or_tmp)
      | (CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0!=5'b00000) | and_830_cse |
      mux_tmp_472);
  assign nor_301_nl = ~(lfst_exit_STORE_LOOP_lpi_2_1 | lfst_exit_STORE_LOOP_lpi_2_0
      | (~ lfst_exit_STORE_LOOP_lpi_2_2) | (CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0!=5'b00000)
      | exitL_exit_STORE_LOOP_sva | mux_tmp_472);
  assign mux_498_nl = MUX_s_1_2_2(nor_300_nl, nor_301_nl, or_214_cse);
  assign CONVOLUTION_LOOP_for_for_for_if_and_cse = core_wen & ((mux_498_nl & BATCH_LOOP_and_6_tmp
      & (fsm_output[2])) | or_tmp_805);
  assign nor_296_nl = ~(lfst_exit_STORE_LOOP_lpi_2_0 | (~(BATCH_LOOP_stage_0 | BATCH_LOOP_stage_0_1
      | BATCH_LOOP_stage_0_3 | BATCH_LOOP_stage_0_4 | (~ or_tmp_16))));
  assign nor_298_nl = ~(STORE_LOOP_or_2336_tmp | not_tmp_291);
  assign nor_299_nl = ~(lfst_exit_STORE_LOOP_lpi_2_0 | not_tmp_291);
  assign mux_514_nl = MUX_s_1_2_2(nor_298_nl, nor_299_nl, BATCH_LOOP_asn_itm_1);
  assign mux_515_nl = MUX_s_1_2_2(nor_296_nl, mux_514_nl, BATCH_LOOP_and_4_tmp);
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_11_cse = core_wen & mux_515_nl & BATCH_LOOP_and_6_tmp
      & (fsm_output[2]);
  assign or_306_cse = (~((~ BATCH_LOOP_if_2_equal_tmp) | (operator_8_false_11_acc_tmp[8:4]!=5'b00000)))
      | (BATCH_LOOP_acc_1_tmp[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_837_cse = core_wen & (~((~ (fsm_output[2]))
      | (and_dcpl_109 & and_dcpl_107) | or_dcpl_51 | (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse)
      | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse | (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1)));
  assign nor_253_nl = ~(nor_303_cse | STORE_LOOP_or_2336_tmp | mux_tmp_512);
  assign nor_255_nl = ~(nor_306_cse | lfst_exit_STORE_LOOP_lpi_2_0 | mux_tmp_510);
  assign mux_520_nl = MUX_s_1_2_2(nor_253_nl, nor_255_nl, or_214_cse);
  assign CONVOLUTION_LOOP_for_for_for_else_and_841_cse = core_wen & (fsm_output[2])
      & mux_520_nl & BATCH_LOOP_and_6_tmp;
  assign nor_249_nl = ~((CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0!=5'b00000)
      | STORE_LOOP_or_2336_tmp | mux_tmp_512);
  assign nor_250_nl = ~((CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0!=5'b00000) | lfst_exit_STORE_LOOP_lpi_2_0
      | mux_tmp_510);
  assign mux_524_nl = MUX_s_1_2_2(nor_249_nl, nor_250_nl, or_214_cse);
  assign CONVOLUTION_LOOP_for_for_for_if_and_833_cse = core_wen & (fsm_output[2])
      & mux_524_nl & BATCH_LOOP_and_6_tmp;
  assign CONVOLUTION_LOOP_for_for_and_3_cse = core_wen & (((~ mux_tmp_468) & BATCH_LOOP_and_6_tmp
      & (fsm_output[2])) | or_tmp_841);
  assign CONVOLUTION_LOOP_for_for_for_acc_and_1_cse = core_wen & ((mux_tmp_351 &
      and_dcpl_22 & STORE_LOOP_equal_tmp_2_2 & (fsm_output[2])) | or_tmp_851);
  assign dma_read_info_index_and_itm = core_wen & BATCH_LOOP_and_6_tmp;
  assign STORE_LOOP_and_726_cse = core_wen & BATCH_LOOP_and_4_tmp;
  assign and_986_cse = core_wen & (~ (fsm_output[2]));
  assign PADDING_LOOP_for_row_and_1_rgt = (~ or_dcpl_60) & (fsm_output[2]);
  assign PADDING_LOOP_for_row_and_3_cse = core_wen & ((~ (fsm_output[2])) | PADDING_LOOP_for_row_and_1_rgt);
  assign PADDING_LOOP_for_and_3_cse = core_wen & (~(or_dcpl_60 & (fsm_output[2])));
  assign or_141_cse = lfst_exit_STORE_LOOP_lpi_2_1 | (~ lfst_exit_STORE_LOOP_lpi_2_2)
      | exitL_exit_STORE_LOOP_sva;
  assign CONVOLUTION_LOOP_for_for_for_for_and_12_cse = core_wen & (~(or_dcpl_85 &
      (fsm_output[2])));
  assign CONVOLUTION_LOOP_for_for_for_y_and_4_rgt = (~ or_dcpl_85) & (fsm_output[2]);
  assign CONVOLUTION_LOOP_for_for_for_y_and_2_rgt = (~(or_tmp_645 | (~ BATCH_LOOP_and_6_tmp)))
      & (fsm_output[2]);
  assign or_1123_tmp = or_dcpl_135 | STORE_LOOP_equal_tmp_4 | STORE_LOOP_equal_tmp_2_mx0w0
      | (STORE_LOOP_equal_tmp_5 & (~ PADDING_LOOP_for_and_tmp_1)) | STORE_LOOP_and_29_cse;
  assign STORE_LOOP_and_22_tmp = PADDING_LOOP_for_and_tmp_1 & STORE_LOOP_equal_tmp_5;
  assign nor_388_nl = ~(STORE_LOOP_and_22_tmp | or_1123_tmp);
  assign PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0_mx1w0 = MUX1HOT_v_5_3_2((signext_5_1(~
      exit_LOAD_LOOP_lpi_2_dfm_1)), (PADDING_LOOP_chan_5_0_sva_2[4:0]), PADDING_LOOP_chan_5_0_lpi_2_4_0,
      {nor_388_nl , STORE_LOOP_and_22_tmp , or_1123_tmp});
  assign exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0 = (~ operator_8_false_2_acc_itm_4_1)
      | exit_PADDING_LOOP_for_sva_5;
  assign exit_CONVOLUTION_LOOP_lpi_2_dfm_mx0w0 = (CONVOLUTION_LOOP_acc_tmp[5]) |
      exit_CONVOLUTION_LOOP_sva_2;
  assign or_1127_tmp = or_dcpl_135 | STORE_LOOP_and_31_cse | (STORE_LOOP_equal_tmp_2_mx0w0
      & (~ CONVOLUTION_LOOP_for_and_tmp_1)) | STORE_LOOP_equal_tmp_4 | STORE_LOOP_equal_tmp_6;
  assign STORE_LOOP_and_24_tmp = CONVOLUTION_LOOP_for_and_tmp_1 & STORE_LOOP_equal_tmp_2_mx0w0;
  assign nor_389_nl = ~(STORE_LOOP_and_24_tmp | or_1127_tmp);
  assign CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0_mx1w0 = MUX1HOT_v_5_3_2((signext_5_1(~
      exit_PADDING_LOOP_lpi_2_dfm_3)), (CONVOLUTION_LOOP_acc_tmp[4:0]), CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0,
      {nor_389_nl , STORE_LOOP_and_24_tmp , or_1127_tmp});
  assign exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0 = (CONVOLUTION_LOOP_for_acc_tmp[5])
      | CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_mx0w0;
  assign exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0 = ~(operator_8_false_6_acc_itm_4_1
      & ((~(CONVOLUTION_LOOP_for_for_if_equal_tmp & (operator_8_false_8_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_8_acc_tmp[8])));
  assign exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1_mx0w0 = (~ operator_8_false_8_acc_itm_3_1)
      | exit_CONVOLUTION_LOOP_for_for_for_for_sva_5;
  assign lfst_exit_STORE_LOOP_lpi_2_2_mx1 = MUX_s_1_2_2(STORE_LOOP_STORE_LOOP_or_tmp,
      lfst_exit_STORE_LOOP_lpi_2_2, or_214_cse);
  assign lfst_exit_STORE_LOOP_lpi_2_0_mx1 = MUX_s_1_2_2(STORE_LOOP_or_2336_tmp, lfst_exit_STORE_LOOP_lpi_2_0,
      or_214_cse);
  assign lfst_exit_STORE_LOOP_lpi_2_1_mx1 = MUX_s_1_2_2(STORE_LOOP_or_2335_tmp, lfst_exit_STORE_LOOP_lpi_2_1,
      or_214_cse);
  assign PADDING_LOOP_for_for_land_2_lpi_2_dfm_mx1w0 = (z_out_2[9]) & PADDING_LOOP_for_for_aelse_1_acc_itm_9_1
      & (~((z_out_1_8_0[8]) | (z_out_3[8])));
  assign exit_BATCH_LOOP_lpi_2_dfm_2_mx1w0 = ((BATCH_LOOP_acc_1_tmp[4]) | exit_BATCH_LOOP_sva_2)
      & exit_STORE_LOOP_lpi_2_dfm_1 & STORE_LOOP_equal_tmp_4;
  assign CONVOLUTION_LOOP_for_for_mux_3_nl = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_and_psp_mx1w0,
      CONVOLUTION_LOOP_for_for_and_psp, mux_tmp_468);
  assign or_1134_nl = (STORE_LOOP_equal_tmp_2_mx0w0 & exit_CONVOLUTION_LOOP_lpi_2_dfm_mx0w0
      & exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4 & CONVOLUTION_LOOP_for_for_and_psp_mx1w0)
      | (CONVOLUTION_LOOP_for_for_mux_3_nl & (~ exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4)
      & STORE_LOOP_equal_tmp_2_mx0w0);
  assign mux_556_nl = MUX_v_5_2_2(CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1, (CONVOLUTION_LOOP_for_acc_tmp[4:0]),
      or_1134_nl);
  assign nor_399_nl = ~((STORE_LOOP_equal_tmp_2_mx0w0 & (~ exit_CONVOLUTION_LOOP_lpi_2_dfm_mx0w0)
      & exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4) | STORE_LOOP_and_32_cse);
  assign CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0_mx1w0 = MUX_v_5_2_2(5'b00000,
      mux_556_nl, nor_399_nl);
  assign lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0 = lfst_exit_STORE_LOOP_lpi_2_2_mx1
      & (~ exitL_exit_STORE_LOOP_sva_mx1);
  assign STORE_LOOP_or_tmp_mx0w0 = (lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1 & (~(lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0
      | lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1))) | (~(lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0
      | lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1 | lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1));
  assign lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1 = lfst_exit_STORE_LOOP_lpi_2_0_mx1
      & (~ exitL_exit_STORE_LOOP_sva_mx1);
  assign lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1 = lfst_exit_STORE_LOOP_lpi_2_1_mx1
      & (~ exitL_exit_STORE_LOOP_sva_mx1);
  assign or_474_nl = (z_out_4[7:6]!=2'b00) | (~ CONVOLUTION_LOOP_for_for_for_if_1_equal_cse)
      | (z_out_4[5]) | (z_out_4[8]) | or_tmp_405;
  assign mux_369_nl = MUX_s_1_2_2(or_474_nl, or_tmp_405, CONVOLUTION_LOOP_for_acc_tmp[5]);
  assign or_475_nl = and_769_cse | mux_369_nl;
  assign CONVOLUTION_LOOP_mux_1_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_lpi_2_dfm_mx0w0,
      exit_CONVOLUTION_LOOP_lpi_2_dfm, or_475_nl);
  assign exit_CONVOLUTION_LOOP_lpi_2_dfm_2_mx0w0 = CONVOLUTION_LOOP_mux_1_nl & exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4;
  assign STORE_LOOP_equal_tmp_2_mx0w0 = lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0 &
      (~(lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1 | lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1));
  assign CONVOLUTION_LOOP_for_for_for_if_1_equal_cse = CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1
      == (z_out_4[4:0]);
  assign CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_mx0w0
      = ~((~(CONVOLUTION_LOOP_for_for_for_if_1_equal_cse & CONVOLUTION_LOOP_for_if_nor_cse))
      | (z_out_4[8]));
  assign PADDING_LOOP_for_for_and_psp_mx1w0 = (~ exit_PADDING_LOOP_for_sva_5) & exit_PADDING_LOOP_for_for_lpi_2_dfm_1;
  assign exit_PADDING_LOOP_lpi_2_dfm_mx0w0 = (PADDING_LOOP_chan_5_0_sva_2[5]) | exit_PADDING_LOOP_sva_2;
  assign CONVOLUTION_LOOP_for_for_and_psp_mx1w0 = (~ CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_mx0w0)
      & exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4;
  assign CONVOLUTION_LOOP_for_for_for_acc_and_4_nl = STORE_LOOP_equal_tmp_2_2 & (~
      or_dcpl_88);
  assign CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_mx1 = MUX_v_45_2_2(CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, CONVOLUTION_LOOP_for_for_for_acc_and_4_nl);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_mx0w0 = MUX_s_1_324_2(buf_acc_data_0_0_0_sva_mx0,
      buf_acc_data_0_1_0_sva_mx0, buf_acc_data_0_2_0_sva_mx0, buf_acc_data_0_3_0_sva_mx0,
      buf_acc_data_0_4_0_sva_mx0, buf_acc_data_0_5_0_sva_mx0, buf_acc_data_0_6_0_sva_mx0,
      buf_acc_data_0_7_0_sva_mx0, buf_acc_data_0_8_0_sva_mx0, buf_acc_data_0_9_0_sva_mx0,
      buf_acc_data_0_10_0_sva_mx0, buf_acc_data_0_11_0_sva_mx0, buf_acc_data_0_12_0_sva_mx0,
      buf_acc_data_0_13_0_sva_mx0, buf_acc_data_0_14_0_sva_mx0, buf_acc_data_0_15_0_sva_mx0,
      buf_acc_data_0_16_0_sva_mx0, buf_acc_data_0_17_0_sva_mx0, buf_acc_data_1_0_0_sva_mx0,
      buf_acc_data_1_1_0_sva_mx0, buf_acc_data_1_2_0_sva_mx0, buf_acc_data_1_3_0_sva_mx0,
      buf_acc_data_1_4_0_sva_mx0, buf_acc_data_1_5_0_sva_mx0, buf_acc_data_1_6_0_sva_mx0,
      buf_acc_data_1_7_0_sva_mx0, buf_acc_data_1_8_0_sva_mx0, buf_acc_data_1_9_0_sva_mx0,
      buf_acc_data_1_10_0_sva_mx0, buf_acc_data_1_11_0_sva_mx0, buf_acc_data_1_12_0_sva_mx0,
      buf_acc_data_1_13_0_sva_mx0, buf_acc_data_1_14_0_sva_mx0, buf_acc_data_1_15_0_sva_mx0,
      buf_acc_data_1_16_0_sva_mx0, buf_acc_data_1_17_0_sva_mx0, buf_acc_data_2_0_0_sva_mx0,
      buf_acc_data_2_1_0_sva_mx0, buf_acc_data_2_2_0_sva_mx0, buf_acc_data_2_3_0_sva_mx0,
      buf_acc_data_2_4_0_sva_mx0, buf_acc_data_2_5_0_sva_mx0, buf_acc_data_2_6_0_sva_mx0,
      buf_acc_data_2_7_0_sva_mx0, buf_acc_data_2_8_0_sva_mx0, buf_acc_data_2_9_0_sva_mx0,
      buf_acc_data_2_10_0_sva_mx0, buf_acc_data_2_11_0_sva_mx0, buf_acc_data_2_12_0_sva_mx0,
      buf_acc_data_2_13_0_sva_mx0, buf_acc_data_2_14_0_sva_mx0, buf_acc_data_2_15_0_sva_mx0,
      buf_acc_data_2_16_0_sva_mx0, buf_acc_data_2_17_0_sva_mx0, buf_acc_data_3_0_0_sva_mx0,
      buf_acc_data_3_1_0_sva_mx0, buf_acc_data_3_2_0_sva_mx0, buf_acc_data_3_3_0_sva_mx0,
      buf_acc_data_3_4_0_sva_mx0, buf_acc_data_3_5_0_sva_mx0, buf_acc_data_3_6_0_sva_mx0,
      buf_acc_data_3_7_0_sva_mx0, buf_acc_data_3_8_0_sva_mx0, buf_acc_data_3_9_0_sva_mx0,
      buf_acc_data_3_10_0_sva_mx0, buf_acc_data_3_11_0_sva_mx0, buf_acc_data_3_12_0_sva_mx0,
      buf_acc_data_3_13_0_sva_mx0, buf_acc_data_3_14_0_sva_mx0, buf_acc_data_3_15_0_sva_mx0,
      buf_acc_data_3_16_0_sva_mx0, buf_acc_data_3_17_0_sva_mx0, buf_acc_data_4_0_0_sva_mx0,
      buf_acc_data_4_1_0_sva_mx0, buf_acc_data_4_2_0_sva_mx0, buf_acc_data_4_3_0_sva_mx0,
      buf_acc_data_4_4_0_sva_mx0, buf_acc_data_4_5_0_sva_mx0, buf_acc_data_4_6_0_sva_mx0,
      buf_acc_data_4_7_0_sva_mx0, buf_acc_data_4_8_0_sva_mx0, buf_acc_data_4_9_0_sva_mx0,
      buf_acc_data_4_10_0_sva_mx0, buf_acc_data_4_11_0_sva_mx0, buf_acc_data_4_12_0_sva_mx0,
      buf_acc_data_4_13_0_sva_mx0, buf_acc_data_4_14_0_sva_mx0, buf_acc_data_4_15_0_sva_mx0,
      buf_acc_data_4_16_0_sva_mx0, buf_acc_data_4_17_0_sva_mx0, buf_acc_data_5_0_0_sva_mx0,
      buf_acc_data_5_1_0_sva_mx0, buf_acc_data_5_2_0_sva_mx0, buf_acc_data_5_3_0_sva_mx0,
      buf_acc_data_5_4_0_sva_mx0, buf_acc_data_5_5_0_sva_mx0, buf_acc_data_5_6_0_sva_mx0,
      buf_acc_data_5_7_0_sva_mx0, buf_acc_data_5_8_0_sva_mx0, buf_acc_data_5_9_0_sva_mx0,
      buf_acc_data_5_10_0_sva_mx0, buf_acc_data_5_11_0_sva_mx0, buf_acc_data_5_12_0_sva_mx0,
      buf_acc_data_5_13_0_sva_mx0, buf_acc_data_5_14_0_sva_mx0, buf_acc_data_5_15_0_sva_mx0,
      buf_acc_data_5_16_0_sva_mx0, buf_acc_data_5_17_0_sva_mx0, buf_acc_data_6_0_0_sva_mx0,
      buf_acc_data_6_1_0_sva_mx0, buf_acc_data_6_2_0_sva_mx0, buf_acc_data_6_3_0_sva_mx0,
      buf_acc_data_6_4_0_sva_mx0, buf_acc_data_6_5_0_sva_mx0, buf_acc_data_6_6_0_sva_mx0,
      buf_acc_data_6_7_0_sva_mx0, buf_acc_data_6_8_0_sva_mx0, buf_acc_data_6_9_0_sva_mx0,
      buf_acc_data_6_10_0_sva_mx0, buf_acc_data_6_11_0_sva_mx0, buf_acc_data_6_12_0_sva_mx0,
      buf_acc_data_6_13_0_sva_mx0, buf_acc_data_6_14_0_sva_mx0, buf_acc_data_6_15_0_sva_mx0,
      buf_acc_data_6_16_0_sva_mx0, buf_acc_data_6_17_0_sva_mx0, buf_acc_data_7_0_0_sva_mx0,
      buf_acc_data_7_1_0_sva_mx0, buf_acc_data_7_2_0_sva_mx0, buf_acc_data_7_3_0_sva_mx0,
      buf_acc_data_7_4_0_sva_mx0, buf_acc_data_7_5_0_sva_mx0, buf_acc_data_7_6_0_sva_mx0,
      buf_acc_data_7_7_0_sva_mx0, buf_acc_data_7_8_0_sva_mx0, buf_acc_data_7_9_0_sva_mx0,
      buf_acc_data_7_10_0_sva_mx0, buf_acc_data_7_11_0_sva_mx0, buf_acc_data_7_12_0_sva_mx0,
      buf_acc_data_7_13_0_sva_mx0, buf_acc_data_7_14_0_sva_mx0, buf_acc_data_7_15_0_sva_mx0,
      buf_acc_data_7_16_0_sva_mx0, buf_acc_data_7_17_0_sva_mx0, buf_acc_data_8_0_0_sva_mx0,
      buf_acc_data_8_1_0_sva_mx0, buf_acc_data_8_2_0_sva_mx0, buf_acc_data_8_3_0_sva_mx0,
      buf_acc_data_8_4_0_sva_mx0, buf_acc_data_8_5_0_sva_mx0, buf_acc_data_8_6_0_sva_mx0,
      buf_acc_data_8_7_0_sva_mx0, buf_acc_data_8_8_0_sva_mx0, buf_acc_data_8_9_0_sva_mx0,
      buf_acc_data_8_10_0_sva_mx0, buf_acc_data_8_11_0_sva_mx0, buf_acc_data_8_12_0_sva_mx0,
      buf_acc_data_8_13_0_sva_mx0, buf_acc_data_8_14_0_sva_mx0, buf_acc_data_8_15_0_sva_mx0,
      buf_acc_data_8_16_0_sva_mx0, buf_acc_data_8_17_0_sva_mx0, buf_acc_data_9_0_0_sva_mx0,
      buf_acc_data_9_1_0_sva_mx0, buf_acc_data_9_2_0_sva_mx0, buf_acc_data_9_3_0_sva_mx0,
      buf_acc_data_9_4_0_sva_mx0, buf_acc_data_9_5_0_sva_mx0, buf_acc_data_9_6_0_sva_mx0,
      buf_acc_data_9_7_0_sva_mx0, buf_acc_data_9_8_0_sva_mx0, buf_acc_data_9_9_0_sva_mx0,
      buf_acc_data_9_10_0_sva_mx0, buf_acc_data_9_11_0_sva_mx0, buf_acc_data_9_12_0_sva_mx0,
      buf_acc_data_9_13_0_sva_mx0, buf_acc_data_9_14_0_sva_mx0, buf_acc_data_9_15_0_sva_mx0,
      buf_acc_data_9_16_0_sva_mx0, buf_acc_data_9_17_0_sva_mx0, buf_acc_data_10_0_0_sva_mx0,
      buf_acc_data_10_1_0_sva_mx0, buf_acc_data_10_2_0_sva_mx0, buf_acc_data_10_3_0_sva_mx0,
      buf_acc_data_10_4_0_sva_mx0, buf_acc_data_10_5_0_sva_mx0, buf_acc_data_10_6_0_sva_mx0,
      buf_acc_data_10_7_0_sva_mx0, buf_acc_data_10_8_0_sva_mx0, buf_acc_data_10_9_0_sva_mx0,
      buf_acc_data_10_10_0_sva_mx0, buf_acc_data_10_11_0_sva_mx0, buf_acc_data_10_12_0_sva_mx0,
      buf_acc_data_10_13_0_sva_mx0, buf_acc_data_10_14_0_sva_mx0, buf_acc_data_10_15_0_sva_mx0,
      buf_acc_data_10_16_0_sva_mx0, buf_acc_data_10_17_0_sva_mx0, buf_acc_data_11_0_0_sva_mx0,
      buf_acc_data_11_1_0_sva_mx0, buf_acc_data_11_2_0_sva_mx0, buf_acc_data_11_3_0_sva_mx0,
      buf_acc_data_11_4_0_sva_mx0, buf_acc_data_11_5_0_sva_mx0, buf_acc_data_11_6_0_sva_mx0,
      buf_acc_data_11_7_0_sva_mx0, buf_acc_data_11_8_0_sva_mx0, buf_acc_data_11_9_0_sva_mx0,
      buf_acc_data_11_10_0_sva_mx0, buf_acc_data_11_11_0_sva_mx0, buf_acc_data_11_12_0_sva_mx0,
      buf_acc_data_11_13_0_sva_mx0, buf_acc_data_11_14_0_sva_mx0, buf_acc_data_11_15_0_sva_mx0,
      buf_acc_data_11_16_0_sva_mx0, buf_acc_data_11_17_0_sva_mx0, buf_acc_data_12_0_0_sva_mx0,
      buf_acc_data_12_1_0_sva_mx0, buf_acc_data_12_2_0_sva_mx0, buf_acc_data_12_3_0_sva_mx0,
      buf_acc_data_12_4_0_sva_mx0, buf_acc_data_12_5_0_sva_mx0, buf_acc_data_12_6_0_sva_mx0,
      buf_acc_data_12_7_0_sva_mx0, buf_acc_data_12_8_0_sva_mx0, buf_acc_data_12_9_0_sva_mx0,
      buf_acc_data_12_10_0_sva_mx0, buf_acc_data_12_11_0_sva_mx0, buf_acc_data_12_12_0_sva_mx0,
      buf_acc_data_12_13_0_sva_mx0, buf_acc_data_12_14_0_sva_mx0, buf_acc_data_12_15_0_sva_mx0,
      buf_acc_data_12_16_0_sva_mx0, buf_acc_data_12_17_0_sva_mx0, buf_acc_data_13_0_0_sva_mx0,
      buf_acc_data_13_1_0_sva_mx0, buf_acc_data_13_2_0_sva_mx0, buf_acc_data_13_3_0_sva_mx0,
      buf_acc_data_13_4_0_sva_mx0, buf_acc_data_13_5_0_sva_mx0, buf_acc_data_13_6_0_sva_mx0,
      buf_acc_data_13_7_0_sva_mx0, buf_acc_data_13_8_0_sva_mx0, buf_acc_data_13_9_0_sva_mx0,
      buf_acc_data_13_10_0_sva_mx0, buf_acc_data_13_11_0_sva_mx0, buf_acc_data_13_12_0_sva_mx0,
      buf_acc_data_13_13_0_sva_mx0, buf_acc_data_13_14_0_sva_mx0, buf_acc_data_13_15_0_sva_mx0,
      buf_acc_data_13_16_0_sva_mx0, buf_acc_data_13_17_0_sva_mx0, buf_acc_data_14_0_0_sva_mx0,
      buf_acc_data_14_1_0_sva_mx0, buf_acc_data_14_2_0_sva_mx0, buf_acc_data_14_3_0_sva_mx0,
      buf_acc_data_14_4_0_sva_mx0, buf_acc_data_14_5_0_sva_mx0, buf_acc_data_14_6_0_sva_mx0,
      buf_acc_data_14_7_0_sva_mx0, buf_acc_data_14_8_0_sva_mx0, buf_acc_data_14_9_0_sva_mx0,
      buf_acc_data_14_10_0_sva_mx0, buf_acc_data_14_11_0_sva_mx0, buf_acc_data_14_12_0_sva_mx0,
      buf_acc_data_14_13_0_sva_mx0, buf_acc_data_14_14_0_sva_mx0, buf_acc_data_14_15_0_sva_mx0,
      buf_acc_data_14_16_0_sva_mx0, buf_acc_data_14_17_0_sva_mx0, buf_acc_data_15_0_0_sva_mx0,
      buf_acc_data_15_1_0_sva_mx0, buf_acc_data_15_2_0_sva_mx0, buf_acc_data_15_3_0_sva_mx0,
      buf_acc_data_15_4_0_sva_mx0, buf_acc_data_15_5_0_sva_mx0, buf_acc_data_15_6_0_sva_mx0,
      buf_acc_data_15_7_0_sva_mx0, buf_acc_data_15_8_0_sva_mx0, buf_acc_data_15_9_0_sva_mx0,
      buf_acc_data_15_10_0_sva_mx0, buf_acc_data_15_11_0_sva_mx0, buf_acc_data_15_12_0_sva_mx0,
      buf_acc_data_15_13_0_sva_mx0, buf_acc_data_15_14_0_sva_mx0, buf_acc_data_15_15_0_sva_mx0,
      buf_acc_data_15_16_0_sva_mx0, buf_acc_data_15_17_0_sva_mx0, buf_acc_data_16_0_0_sva_mx0,
      buf_acc_data_16_1_0_sva_mx0, buf_acc_data_16_2_0_sva_mx0, buf_acc_data_16_3_0_sva_mx0,
      buf_acc_data_16_4_0_sva_mx0, buf_acc_data_16_5_0_sva_mx0, buf_acc_data_16_6_0_sva_mx0,
      buf_acc_data_16_7_0_sva_mx0, buf_acc_data_16_8_0_sva_mx0, buf_acc_data_16_9_0_sva_mx0,
      buf_acc_data_16_10_0_sva_mx0, buf_acc_data_16_11_0_sva_mx0, buf_acc_data_16_12_0_sva_mx0,
      buf_acc_data_16_13_0_sva_mx0, buf_acc_data_16_14_0_sva_mx0, buf_acc_data_16_15_0_sva_mx0,
      buf_acc_data_16_16_0_sva_mx0, buf_acc_data_16_17_0_sva_mx0, buf_acc_data_17_0_0_sva_mx0,
      buf_acc_data_17_1_0_sva_mx0, buf_acc_data_17_2_0_sva_mx0, buf_acc_data_17_3_0_sva_mx0,
      buf_acc_data_17_4_0_sva_mx0, buf_acc_data_17_5_0_sva_mx0, buf_acc_data_17_6_0_sva_mx0,
      buf_acc_data_17_7_0_sva_mx0, buf_acc_data_17_8_0_sva_mx0, buf_acc_data_17_9_0_sva_mx0,
      buf_acc_data_17_10_0_sva_mx0, buf_acc_data_17_11_0_sva_mx0, buf_acc_data_17_12_0_sva_mx0,
      buf_acc_data_17_13_0_sva_mx0, buf_acc_data_17_14_0_sva_mx0, buf_acc_data_17_15_0_sva_mx0,
      buf_acc_data_17_16_0_sva_mx0, buf_acc_data_17_17_0_sva_mx0, {CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3
      , CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_1_0});
  assign CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_mx0w0 = MUX_v_45_324_2(buf_acc_data_0_0_45_1_sva_mx0,
      buf_acc_data_0_1_45_1_sva_mx0, buf_acc_data_0_2_45_1_sva_mx0, buf_acc_data_0_3_45_1_sva_mx0,
      buf_acc_data_0_4_45_1_sva_mx0, buf_acc_data_0_5_45_1_sva_mx0, buf_acc_data_0_6_45_1_sva_mx0,
      buf_acc_data_0_7_45_1_sva_mx0, buf_acc_data_0_8_45_1_sva_mx0, buf_acc_data_0_9_45_1_sva_mx0,
      buf_acc_data_0_10_45_1_sva_mx0, buf_acc_data_0_11_45_1_sva_mx0, buf_acc_data_0_12_45_1_sva_mx0,
      buf_acc_data_0_13_45_1_sva_mx0, buf_acc_data_0_14_45_1_sva_mx0, buf_acc_data_0_15_45_1_sva_mx0,
      buf_acc_data_0_16_45_1_sva_mx0, buf_acc_data_0_17_45_1_sva_mx0, buf_acc_data_1_0_45_1_sva_mx0,
      buf_acc_data_1_1_45_1_sva_mx0, buf_acc_data_1_2_45_1_sva_mx0, buf_acc_data_1_3_45_1_sva_mx0,
      buf_acc_data_1_4_45_1_sva_mx0, buf_acc_data_1_5_45_1_sva_mx0, buf_acc_data_1_6_45_1_sva_mx0,
      buf_acc_data_1_7_45_1_sva_mx0, buf_acc_data_1_8_45_1_sva_mx0, buf_acc_data_1_9_45_1_sva_mx0,
      buf_acc_data_1_10_45_1_sva_mx0, buf_acc_data_1_11_45_1_sva_mx0, buf_acc_data_1_12_45_1_sva_mx0,
      buf_acc_data_1_13_45_1_sva_mx0, buf_acc_data_1_14_45_1_sva_mx0, buf_acc_data_1_15_45_1_sva_mx0,
      buf_acc_data_1_16_45_1_sva_mx0, buf_acc_data_1_17_45_1_sva_mx0, buf_acc_data_2_0_45_1_sva_mx0,
      buf_acc_data_2_1_45_1_sva_mx0, buf_acc_data_2_2_45_1_sva_mx0, buf_acc_data_2_3_45_1_sva_mx0,
      buf_acc_data_2_4_45_1_sva_mx0, buf_acc_data_2_5_45_1_sva_mx0, buf_acc_data_2_6_45_1_sva_mx0,
      buf_acc_data_2_7_45_1_sva_mx0, buf_acc_data_2_8_45_1_sva_mx0, buf_acc_data_2_9_45_1_sva_mx0,
      buf_acc_data_2_10_45_1_sva_mx0, buf_acc_data_2_11_45_1_sva_mx0, buf_acc_data_2_12_45_1_sva_mx0,
      buf_acc_data_2_13_45_1_sva_mx0, buf_acc_data_2_14_45_1_sva_mx0, buf_acc_data_2_15_45_1_sva_mx0,
      buf_acc_data_2_16_45_1_sva_mx0, buf_acc_data_2_17_45_1_sva_mx0, buf_acc_data_3_0_45_1_sva_mx0,
      buf_acc_data_3_1_45_1_sva_mx0, buf_acc_data_3_2_45_1_sva_mx0, buf_acc_data_3_3_45_1_sva_mx0,
      buf_acc_data_3_4_45_1_sva_mx0, buf_acc_data_3_5_45_1_sva_mx0, buf_acc_data_3_6_45_1_sva_mx0,
      buf_acc_data_3_7_45_1_sva_mx0, buf_acc_data_3_8_45_1_sva_mx0, buf_acc_data_3_9_45_1_sva_mx0,
      buf_acc_data_3_10_45_1_sva_mx0, buf_acc_data_3_11_45_1_sva_mx0, buf_acc_data_3_12_45_1_sva_mx0,
      buf_acc_data_3_13_45_1_sva_mx0, buf_acc_data_3_14_45_1_sva_mx0, buf_acc_data_3_15_45_1_sva_mx0,
      buf_acc_data_3_16_45_1_sva_mx0, buf_acc_data_3_17_45_1_sva_mx0, buf_acc_data_4_0_45_1_sva_mx0,
      buf_acc_data_4_1_45_1_sva_mx0, buf_acc_data_4_2_45_1_sva_mx0, buf_acc_data_4_3_45_1_sva_mx0,
      buf_acc_data_4_4_45_1_sva_mx0, buf_acc_data_4_5_45_1_sva_mx0, buf_acc_data_4_6_45_1_sva_mx0,
      buf_acc_data_4_7_45_1_sva_mx0, buf_acc_data_4_8_45_1_sva_mx0, buf_acc_data_4_9_45_1_sva_mx0,
      buf_acc_data_4_10_45_1_sva_mx0, buf_acc_data_4_11_45_1_sva_mx0, buf_acc_data_4_12_45_1_sva_mx0,
      buf_acc_data_4_13_45_1_sva_mx0, buf_acc_data_4_14_45_1_sva_mx0, buf_acc_data_4_15_45_1_sva_mx0,
      buf_acc_data_4_16_45_1_sva_mx0, buf_acc_data_4_17_45_1_sva_mx0, buf_acc_data_5_0_45_1_sva_mx0,
      buf_acc_data_5_1_45_1_sva_mx0, buf_acc_data_5_2_45_1_sva_mx0, buf_acc_data_5_3_45_1_sva_mx0,
      buf_acc_data_5_4_45_1_sva_mx0, buf_acc_data_5_5_45_1_sva_mx0, buf_acc_data_5_6_45_1_sva_mx0,
      buf_acc_data_5_7_45_1_sva_mx0, buf_acc_data_5_8_45_1_sva_mx0, buf_acc_data_5_9_45_1_sva_mx0,
      buf_acc_data_5_10_45_1_sva_mx0, buf_acc_data_5_11_45_1_sva_mx0, buf_acc_data_5_12_45_1_sva_mx0,
      buf_acc_data_5_13_45_1_sva_mx0, buf_acc_data_5_14_45_1_sva_mx0, buf_acc_data_5_15_45_1_sva_mx0,
      buf_acc_data_5_16_45_1_sva_mx0, buf_acc_data_5_17_45_1_sva_mx0, buf_acc_data_6_0_45_1_sva_mx0,
      buf_acc_data_6_1_45_1_sva_mx0, buf_acc_data_6_2_45_1_sva_mx0, buf_acc_data_6_3_45_1_sva_mx0,
      buf_acc_data_6_4_45_1_sva_mx0, buf_acc_data_6_5_45_1_sva_mx0, buf_acc_data_6_6_45_1_sva_mx0,
      buf_acc_data_6_7_45_1_sva_mx0, buf_acc_data_6_8_45_1_sva_mx0, buf_acc_data_6_9_45_1_sva_mx0,
      buf_acc_data_6_10_45_1_sva_mx0, buf_acc_data_6_11_45_1_sva_mx0, buf_acc_data_6_12_45_1_sva_mx0,
      buf_acc_data_6_13_45_1_sva_mx0, buf_acc_data_6_14_45_1_sva_mx0, buf_acc_data_6_15_45_1_sva_mx0,
      buf_acc_data_6_16_45_1_sva_mx0, buf_acc_data_6_17_45_1_sva_mx0, buf_acc_data_7_0_45_1_sva_mx0,
      buf_acc_data_7_1_45_1_sva_mx0, buf_acc_data_7_2_45_1_sva_mx0, buf_acc_data_7_3_45_1_sva_mx0,
      buf_acc_data_7_4_45_1_sva_mx0, buf_acc_data_7_5_45_1_sva_mx0, buf_acc_data_7_6_45_1_sva_mx0,
      buf_acc_data_7_7_45_1_sva_mx0, buf_acc_data_7_8_45_1_sva_mx0, buf_acc_data_7_9_45_1_sva_mx0,
      buf_acc_data_7_10_45_1_sva_mx0, buf_acc_data_7_11_45_1_sva_mx0, buf_acc_data_7_12_45_1_sva_mx0,
      buf_acc_data_7_13_45_1_sva_mx0, buf_acc_data_7_14_45_1_sva_mx0, buf_acc_data_7_15_45_1_sva_mx0,
      buf_acc_data_7_16_45_1_sva_mx0, buf_acc_data_7_17_45_1_sva_mx0, buf_acc_data_8_0_45_1_sva_mx0,
      buf_acc_data_8_1_45_1_sva_mx0, buf_acc_data_8_2_45_1_sva_mx0, buf_acc_data_8_3_45_1_sva_mx0,
      buf_acc_data_8_4_45_1_sva_mx0, buf_acc_data_8_5_45_1_sva_mx0, buf_acc_data_8_6_45_1_sva_mx0,
      buf_acc_data_8_7_45_1_sva_mx0, buf_acc_data_8_8_45_1_sva_mx0, buf_acc_data_8_9_45_1_sva_mx0,
      buf_acc_data_8_10_45_1_sva_mx0, buf_acc_data_8_11_45_1_sva_mx0, buf_acc_data_8_12_45_1_sva_mx0,
      buf_acc_data_8_13_45_1_sva_mx0, buf_acc_data_8_14_45_1_sva_mx0, buf_acc_data_8_15_45_1_sva_mx0,
      buf_acc_data_8_16_45_1_sva_mx0, buf_acc_data_8_17_45_1_sva_mx0, buf_acc_data_9_0_45_1_sva_mx0,
      buf_acc_data_9_1_45_1_sva_mx0, buf_acc_data_9_2_45_1_sva_mx0, buf_acc_data_9_3_45_1_sva_mx0,
      buf_acc_data_9_4_45_1_sva_mx0, buf_acc_data_9_5_45_1_sva_mx0, buf_acc_data_9_6_45_1_sva_mx0,
      buf_acc_data_9_7_45_1_sva_mx0, buf_acc_data_9_8_45_1_sva_mx0, buf_acc_data_9_9_45_1_sva_mx0,
      buf_acc_data_9_10_45_1_sva_mx0, buf_acc_data_9_11_45_1_sva_mx0, buf_acc_data_9_12_45_1_sva_mx0,
      buf_acc_data_9_13_45_1_sva_mx0, buf_acc_data_9_14_45_1_sva_mx0, buf_acc_data_9_15_45_1_sva_mx0,
      buf_acc_data_9_16_45_1_sva_mx0, buf_acc_data_9_17_45_1_sva_mx0, buf_acc_data_10_0_45_1_sva_mx0,
      buf_acc_data_10_1_45_1_sva_mx0, buf_acc_data_10_2_45_1_sva_mx0, buf_acc_data_10_3_45_1_sva_mx0,
      buf_acc_data_10_4_45_1_sva_mx0, buf_acc_data_10_5_45_1_sva_mx0, buf_acc_data_10_6_45_1_sva_mx0,
      buf_acc_data_10_7_45_1_sva_mx0, buf_acc_data_10_8_45_1_sva_mx0, buf_acc_data_10_9_45_1_sva_mx0,
      buf_acc_data_10_10_45_1_sva_mx0, buf_acc_data_10_11_45_1_sva_mx0, buf_acc_data_10_12_45_1_sva_mx0,
      buf_acc_data_10_13_45_1_sva_mx0, buf_acc_data_10_14_45_1_sva_mx0, buf_acc_data_10_15_45_1_sva_mx0,
      buf_acc_data_10_16_45_1_sva_mx0, buf_acc_data_10_17_45_1_sva_mx0, buf_acc_data_11_0_45_1_sva_mx0,
      buf_acc_data_11_1_45_1_sva_mx0, buf_acc_data_11_2_45_1_sva_mx0, buf_acc_data_11_3_45_1_sva_mx0,
      buf_acc_data_11_4_45_1_sva_mx0, buf_acc_data_11_5_45_1_sva_mx0, buf_acc_data_11_6_45_1_sva_mx0,
      buf_acc_data_11_7_45_1_sva_mx0, buf_acc_data_11_8_45_1_sva_mx0, buf_acc_data_11_9_45_1_sva_mx0,
      buf_acc_data_11_10_45_1_sva_mx0, buf_acc_data_11_11_45_1_sva_mx0, buf_acc_data_11_12_45_1_sva_mx0,
      buf_acc_data_11_13_45_1_sva_mx0, buf_acc_data_11_14_45_1_sva_mx0, buf_acc_data_11_15_45_1_sva_mx0,
      buf_acc_data_11_16_45_1_sva_mx0, buf_acc_data_11_17_45_1_sva_mx0, buf_acc_data_12_0_45_1_sva_mx0,
      buf_acc_data_12_1_45_1_sva_mx0, buf_acc_data_12_2_45_1_sva_mx0, buf_acc_data_12_3_45_1_sva_mx0,
      buf_acc_data_12_4_45_1_sva_mx0, buf_acc_data_12_5_45_1_sva_mx0, buf_acc_data_12_6_45_1_sva_mx0,
      buf_acc_data_12_7_45_1_sva_mx0, buf_acc_data_12_8_45_1_sva_mx0, buf_acc_data_12_9_45_1_sva_mx0,
      buf_acc_data_12_10_45_1_sva_mx0, buf_acc_data_12_11_45_1_sva_mx0, buf_acc_data_12_12_45_1_sva_mx0,
      buf_acc_data_12_13_45_1_sva_mx0, buf_acc_data_12_14_45_1_sva_mx0, buf_acc_data_12_15_45_1_sva_mx0,
      buf_acc_data_12_16_45_1_sva_mx0, buf_acc_data_12_17_45_1_sva_mx0, buf_acc_data_13_0_45_1_sva_mx0,
      buf_acc_data_13_1_45_1_sva_mx0, buf_acc_data_13_2_45_1_sva_mx0, buf_acc_data_13_3_45_1_sva_mx0,
      buf_acc_data_13_4_45_1_sva_mx0, buf_acc_data_13_5_45_1_sva_mx0, buf_acc_data_13_6_45_1_sva_mx0,
      buf_acc_data_13_7_45_1_sva_mx0, buf_acc_data_13_8_45_1_sva_mx0, buf_acc_data_13_9_45_1_sva_mx0,
      buf_acc_data_13_10_45_1_sva_mx0, buf_acc_data_13_11_45_1_sva_mx0, buf_acc_data_13_12_45_1_sva_mx0,
      buf_acc_data_13_13_45_1_sva_mx0, buf_acc_data_13_14_45_1_sva_mx0, buf_acc_data_13_15_45_1_sva_mx0,
      buf_acc_data_13_16_45_1_sva_mx0, buf_acc_data_13_17_45_1_sva_mx0, buf_acc_data_14_0_45_1_sva_mx0,
      buf_acc_data_14_1_45_1_sva_mx0, buf_acc_data_14_2_45_1_sva_mx0, buf_acc_data_14_3_45_1_sva_mx0,
      buf_acc_data_14_4_45_1_sva_mx0, buf_acc_data_14_5_45_1_sva_mx0, buf_acc_data_14_6_45_1_sva_mx0,
      buf_acc_data_14_7_45_1_sva_mx0, buf_acc_data_14_8_45_1_sva_mx0, buf_acc_data_14_9_45_1_sva_mx0,
      buf_acc_data_14_10_45_1_sva_mx0, buf_acc_data_14_11_45_1_sva_mx0, buf_acc_data_14_12_45_1_sva_mx0,
      buf_acc_data_14_13_45_1_sva_mx0, buf_acc_data_14_14_45_1_sva_mx0, buf_acc_data_14_15_45_1_sva_mx0,
      buf_acc_data_14_16_45_1_sva_mx0, buf_acc_data_14_17_45_1_sva_mx0, buf_acc_data_15_0_45_1_sva_mx0,
      buf_acc_data_15_1_45_1_sva_mx0, buf_acc_data_15_2_45_1_sva_mx0, buf_acc_data_15_3_45_1_sva_mx0,
      buf_acc_data_15_4_45_1_sva_mx0, buf_acc_data_15_5_45_1_sva_mx0, buf_acc_data_15_6_45_1_sva_mx0,
      buf_acc_data_15_7_45_1_sva_mx0, buf_acc_data_15_8_45_1_sva_mx0, buf_acc_data_15_9_45_1_sva_mx0,
      buf_acc_data_15_10_45_1_sva_mx0, buf_acc_data_15_11_45_1_sva_mx0, buf_acc_data_15_12_45_1_sva_mx0,
      buf_acc_data_15_13_45_1_sva_mx0, buf_acc_data_15_14_45_1_sva_mx0, buf_acc_data_15_15_45_1_sva_mx0,
      buf_acc_data_15_16_45_1_sva_mx0, buf_acc_data_15_17_45_1_sva_mx0, buf_acc_data_16_0_45_1_sva_mx0,
      buf_acc_data_16_1_45_1_sva_mx0, buf_acc_data_16_2_45_1_sva_mx0, buf_acc_data_16_3_45_1_sva_mx0,
      buf_acc_data_16_4_45_1_sva_mx0, buf_acc_data_16_5_45_1_sva_mx0, buf_acc_data_16_6_45_1_sva_mx0,
      buf_acc_data_16_7_45_1_sva_mx0, buf_acc_data_16_8_45_1_sva_mx0, buf_acc_data_16_9_45_1_sva_mx0,
      buf_acc_data_16_10_45_1_sva_mx0, buf_acc_data_16_11_45_1_sva_mx0, buf_acc_data_16_12_45_1_sva_mx0,
      buf_acc_data_16_13_45_1_sva_mx0, buf_acc_data_16_14_45_1_sva_mx0, buf_acc_data_16_15_45_1_sva_mx0,
      buf_acc_data_16_16_45_1_sva_mx0, buf_acc_data_16_17_45_1_sva_mx0, buf_acc_data_17_0_45_1_sva_mx0,
      buf_acc_data_17_1_45_1_sva_mx0, buf_acc_data_17_2_45_1_sva_mx0, buf_acc_data_17_3_45_1_sva_mx0,
      buf_acc_data_17_4_45_1_sva_mx0, buf_acc_data_17_5_45_1_sva_mx0, buf_acc_data_17_6_45_1_sva_mx0,
      buf_acc_data_17_7_45_1_sva_mx0, buf_acc_data_17_8_45_1_sva_mx0, buf_acc_data_17_9_45_1_sva_mx0,
      buf_acc_data_17_10_45_1_sva_mx0, buf_acc_data_17_11_45_1_sva_mx0, buf_acc_data_17_12_45_1_sva_mx0,
      buf_acc_data_17_13_45_1_sva_mx0, buf_acc_data_17_14_45_1_sva_mx0, buf_acc_data_17_15_45_1_sva_mx0,
      buf_acc_data_17_16_45_1_sva_mx0, buf_acc_data_17_17_45_1_sva_mx0, {CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3
      , CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_1_0});
  assign CONVOLUTION_LOOP_for_for_for_else_mux_itm_mx0w0 = MUX_v_11_324_2(buf_acc_data_0_0_56_46_sva_mx0,
      buf_acc_data_0_1_56_46_sva_mx0, buf_acc_data_0_2_56_46_sva_mx0, buf_acc_data_0_3_56_46_sva_mx0,
      buf_acc_data_0_4_56_46_sva_mx0, buf_acc_data_0_5_56_46_sva_mx0, buf_acc_data_0_6_56_46_sva_mx0,
      buf_acc_data_0_7_56_46_sva_mx0, buf_acc_data_0_8_56_46_sva_mx0, buf_acc_data_0_9_56_46_sva_mx0,
      buf_acc_data_0_10_56_46_sva_mx0, buf_acc_data_0_11_56_46_sva_mx0, buf_acc_data_0_12_56_46_sva_mx0,
      buf_acc_data_0_13_56_46_sva_mx0, buf_acc_data_0_14_56_46_sva_mx0, buf_acc_data_0_15_56_46_sva_mx0,
      buf_acc_data_0_16_56_46_sva_mx0, buf_acc_data_0_17_56_46_sva_mx0, buf_acc_data_1_0_56_46_sva_mx0,
      buf_acc_data_1_1_56_46_sva_mx0, buf_acc_data_1_2_56_46_sva_mx0, buf_acc_data_1_3_56_46_sva_mx0,
      buf_acc_data_1_4_56_46_sva_mx0, buf_acc_data_1_5_56_46_sva_mx0, buf_acc_data_1_6_56_46_sva_mx0,
      buf_acc_data_1_7_56_46_sva_mx0, buf_acc_data_1_8_56_46_sva_mx0, buf_acc_data_1_9_56_46_sva_mx0,
      buf_acc_data_1_10_56_46_sva_mx0, buf_acc_data_1_11_56_46_sva_mx0, buf_acc_data_1_12_56_46_sva_mx0,
      buf_acc_data_1_13_56_46_sva_mx0, buf_acc_data_1_14_56_46_sva_mx0, buf_acc_data_1_15_56_46_sva_mx0,
      buf_acc_data_1_16_56_46_sva_mx0, buf_acc_data_1_17_56_46_sva_mx0, buf_acc_data_2_0_56_46_sva_mx0,
      buf_acc_data_2_1_56_46_sva_mx0, buf_acc_data_2_2_56_46_sva_mx0, buf_acc_data_2_3_56_46_sva_mx0,
      buf_acc_data_2_4_56_46_sva_mx0, buf_acc_data_2_5_56_46_sva_mx0, buf_acc_data_2_6_56_46_sva_mx0,
      buf_acc_data_2_7_56_46_sva_mx0, buf_acc_data_2_8_56_46_sva_mx0, buf_acc_data_2_9_56_46_sva_mx0,
      buf_acc_data_2_10_56_46_sva_mx0, buf_acc_data_2_11_56_46_sva_mx0, buf_acc_data_2_12_56_46_sva_mx0,
      buf_acc_data_2_13_56_46_sva_mx0, buf_acc_data_2_14_56_46_sva_mx0, buf_acc_data_2_15_56_46_sva_mx0,
      buf_acc_data_2_16_56_46_sva_mx0, buf_acc_data_2_17_56_46_sva_mx0, buf_acc_data_3_0_56_46_sva_mx0,
      buf_acc_data_3_1_56_46_sva_mx0, buf_acc_data_3_2_56_46_sva_mx0, buf_acc_data_3_3_56_46_sva_mx0,
      buf_acc_data_3_4_56_46_sva_mx0, buf_acc_data_3_5_56_46_sva_mx0, buf_acc_data_3_6_56_46_sva_mx0,
      buf_acc_data_3_7_56_46_sva_mx0, buf_acc_data_3_8_56_46_sva_mx0, buf_acc_data_3_9_56_46_sva_mx0,
      buf_acc_data_3_10_56_46_sva_mx0, buf_acc_data_3_11_56_46_sva_mx0, buf_acc_data_3_12_56_46_sva_mx0,
      buf_acc_data_3_13_56_46_sva_mx0, buf_acc_data_3_14_56_46_sva_mx0, buf_acc_data_3_15_56_46_sva_mx0,
      buf_acc_data_3_16_56_46_sva_mx0, buf_acc_data_3_17_56_46_sva_mx0, buf_acc_data_4_0_56_46_sva_mx0,
      buf_acc_data_4_1_56_46_sva_mx0, buf_acc_data_4_2_56_46_sva_mx0, buf_acc_data_4_3_56_46_sva_mx0,
      buf_acc_data_4_4_56_46_sva_mx0, buf_acc_data_4_5_56_46_sva_mx0, buf_acc_data_4_6_56_46_sva_mx0,
      buf_acc_data_4_7_56_46_sva_mx0, buf_acc_data_4_8_56_46_sva_mx0, buf_acc_data_4_9_56_46_sva_mx0,
      buf_acc_data_4_10_56_46_sva_mx0, buf_acc_data_4_11_56_46_sva_mx0, buf_acc_data_4_12_56_46_sva_mx0,
      buf_acc_data_4_13_56_46_sva_mx0, buf_acc_data_4_14_56_46_sva_mx0, buf_acc_data_4_15_56_46_sva_mx0,
      buf_acc_data_4_16_56_46_sva_mx0, buf_acc_data_4_17_56_46_sva_mx0, buf_acc_data_5_0_56_46_sva_mx0,
      buf_acc_data_5_1_56_46_sva_mx0, buf_acc_data_5_2_56_46_sva_mx0, buf_acc_data_5_3_56_46_sva_mx0,
      buf_acc_data_5_4_56_46_sva_mx0, buf_acc_data_5_5_56_46_sva_mx0, buf_acc_data_5_6_56_46_sva_mx0,
      buf_acc_data_5_7_56_46_sva_mx0, buf_acc_data_5_8_56_46_sva_mx0, buf_acc_data_5_9_56_46_sva_mx0,
      buf_acc_data_5_10_56_46_sva_mx0, buf_acc_data_5_11_56_46_sva_mx0, buf_acc_data_5_12_56_46_sva_mx0,
      buf_acc_data_5_13_56_46_sva_mx0, buf_acc_data_5_14_56_46_sva_mx0, buf_acc_data_5_15_56_46_sva_mx0,
      buf_acc_data_5_16_56_46_sva_mx0, buf_acc_data_5_17_56_46_sva_mx0, buf_acc_data_6_0_56_46_sva_mx0,
      buf_acc_data_6_1_56_46_sva_mx0, buf_acc_data_6_2_56_46_sva_mx0, buf_acc_data_6_3_56_46_sva_mx0,
      buf_acc_data_6_4_56_46_sva_mx0, buf_acc_data_6_5_56_46_sva_mx0, buf_acc_data_6_6_56_46_sva_mx0,
      buf_acc_data_6_7_56_46_sva_mx0, buf_acc_data_6_8_56_46_sva_mx0, buf_acc_data_6_9_56_46_sva_mx0,
      buf_acc_data_6_10_56_46_sva_mx0, buf_acc_data_6_11_56_46_sva_mx0, buf_acc_data_6_12_56_46_sva_mx0,
      buf_acc_data_6_13_56_46_sva_mx0, buf_acc_data_6_14_56_46_sva_mx0, buf_acc_data_6_15_56_46_sva_mx0,
      buf_acc_data_6_16_56_46_sva_mx0, buf_acc_data_6_17_56_46_sva_mx0, buf_acc_data_7_0_56_46_sva_mx0,
      buf_acc_data_7_1_56_46_sva_mx0, buf_acc_data_7_2_56_46_sva_mx0, buf_acc_data_7_3_56_46_sva_mx0,
      buf_acc_data_7_4_56_46_sva_mx0, buf_acc_data_7_5_56_46_sva_mx0, buf_acc_data_7_6_56_46_sva_mx0,
      buf_acc_data_7_7_56_46_sva_mx0, buf_acc_data_7_8_56_46_sva_mx0, buf_acc_data_7_9_56_46_sva_mx0,
      buf_acc_data_7_10_56_46_sva_mx0, buf_acc_data_7_11_56_46_sva_mx0, buf_acc_data_7_12_56_46_sva_mx0,
      buf_acc_data_7_13_56_46_sva_mx0, buf_acc_data_7_14_56_46_sva_mx0, buf_acc_data_7_15_56_46_sva_mx0,
      buf_acc_data_7_16_56_46_sva_mx0, buf_acc_data_7_17_56_46_sva_mx0, buf_acc_data_8_0_56_46_sva_mx0,
      buf_acc_data_8_1_56_46_sva_mx0, buf_acc_data_8_2_56_46_sva_mx0, buf_acc_data_8_3_56_46_sva_mx0,
      buf_acc_data_8_4_56_46_sva_mx0, buf_acc_data_8_5_56_46_sva_mx0, buf_acc_data_8_6_56_46_sva_mx0,
      buf_acc_data_8_7_56_46_sva_mx0, buf_acc_data_8_8_56_46_sva_mx0, buf_acc_data_8_9_56_46_sva_mx0,
      buf_acc_data_8_10_56_46_sva_mx0, buf_acc_data_8_11_56_46_sva_mx0, buf_acc_data_8_12_56_46_sva_mx0,
      buf_acc_data_8_13_56_46_sva_mx0, buf_acc_data_8_14_56_46_sva_mx0, buf_acc_data_8_15_56_46_sva_mx0,
      buf_acc_data_8_16_56_46_sva_mx0, buf_acc_data_8_17_56_46_sva_mx0, buf_acc_data_9_0_56_46_sva_mx0,
      buf_acc_data_9_1_56_46_sva_mx0, buf_acc_data_9_2_56_46_sva_mx0, buf_acc_data_9_3_56_46_sva_mx0,
      buf_acc_data_9_4_56_46_sva_mx0, buf_acc_data_9_5_56_46_sva_mx0, buf_acc_data_9_6_56_46_sva_mx0,
      buf_acc_data_9_7_56_46_sva_mx0, buf_acc_data_9_8_56_46_sva_mx0, buf_acc_data_9_9_56_46_sva_mx0,
      buf_acc_data_9_10_56_46_sva_mx0, buf_acc_data_9_11_56_46_sva_mx0, buf_acc_data_9_12_56_46_sva_mx0,
      buf_acc_data_9_13_56_46_sva_mx0, buf_acc_data_9_14_56_46_sva_mx0, buf_acc_data_9_15_56_46_sva_mx0,
      buf_acc_data_9_16_56_46_sva_mx0, buf_acc_data_9_17_56_46_sva_mx0, buf_acc_data_10_0_56_46_sva_mx0,
      buf_acc_data_10_1_56_46_sva_mx0, buf_acc_data_10_2_56_46_sva_mx0, buf_acc_data_10_3_56_46_sva_mx0,
      buf_acc_data_10_4_56_46_sva_mx0, buf_acc_data_10_5_56_46_sva_mx0, buf_acc_data_10_6_56_46_sva_mx0,
      buf_acc_data_10_7_56_46_sva_mx0, buf_acc_data_10_8_56_46_sva_mx0, buf_acc_data_10_9_56_46_sva_mx0,
      buf_acc_data_10_10_56_46_sva_mx0, buf_acc_data_10_11_56_46_sva_mx0, buf_acc_data_10_12_56_46_sva_mx0,
      buf_acc_data_10_13_56_46_sva_mx0, buf_acc_data_10_14_56_46_sva_mx0, buf_acc_data_10_15_56_46_sva_mx0,
      buf_acc_data_10_16_56_46_sva_mx0, buf_acc_data_10_17_56_46_sva_mx0, buf_acc_data_11_0_56_46_sva_mx0,
      buf_acc_data_11_1_56_46_sva_mx0, buf_acc_data_11_2_56_46_sva_mx0, buf_acc_data_11_3_56_46_sva_mx0,
      buf_acc_data_11_4_56_46_sva_mx0, buf_acc_data_11_5_56_46_sva_mx0, buf_acc_data_11_6_56_46_sva_mx0,
      buf_acc_data_11_7_56_46_sva_mx0, buf_acc_data_11_8_56_46_sva_mx0, buf_acc_data_11_9_56_46_sva_mx0,
      buf_acc_data_11_10_56_46_sva_mx0, buf_acc_data_11_11_56_46_sva_mx0, buf_acc_data_11_12_56_46_sva_mx0,
      buf_acc_data_11_13_56_46_sva_mx0, buf_acc_data_11_14_56_46_sva_mx0, buf_acc_data_11_15_56_46_sva_mx0,
      buf_acc_data_11_16_56_46_sva_mx0, buf_acc_data_11_17_56_46_sva_mx0, buf_acc_data_12_0_56_46_sva_mx0,
      buf_acc_data_12_1_56_46_sva_mx0, buf_acc_data_12_2_56_46_sva_mx0, buf_acc_data_12_3_56_46_sva_mx0,
      buf_acc_data_12_4_56_46_sva_mx0, buf_acc_data_12_5_56_46_sva_mx0, buf_acc_data_12_6_56_46_sva_mx0,
      buf_acc_data_12_7_56_46_sva_mx0, buf_acc_data_12_8_56_46_sva_mx0, buf_acc_data_12_9_56_46_sva_mx0,
      buf_acc_data_12_10_56_46_sva_mx0, buf_acc_data_12_11_56_46_sva_mx0, buf_acc_data_12_12_56_46_sva_mx0,
      buf_acc_data_12_13_56_46_sva_mx0, buf_acc_data_12_14_56_46_sva_mx0, buf_acc_data_12_15_56_46_sva_mx0,
      buf_acc_data_12_16_56_46_sva_mx0, buf_acc_data_12_17_56_46_sva_mx0, buf_acc_data_13_0_56_46_sva_mx0,
      buf_acc_data_13_1_56_46_sva_mx0, buf_acc_data_13_2_56_46_sva_mx0, buf_acc_data_13_3_56_46_sva_mx0,
      buf_acc_data_13_4_56_46_sva_mx0, buf_acc_data_13_5_56_46_sva_mx0, buf_acc_data_13_6_56_46_sva_mx0,
      buf_acc_data_13_7_56_46_sva_mx0, buf_acc_data_13_8_56_46_sva_mx0, buf_acc_data_13_9_56_46_sva_mx0,
      buf_acc_data_13_10_56_46_sva_mx0, buf_acc_data_13_11_56_46_sva_mx0, buf_acc_data_13_12_56_46_sva_mx0,
      buf_acc_data_13_13_56_46_sva_mx0, buf_acc_data_13_14_56_46_sva_mx0, buf_acc_data_13_15_56_46_sva_mx0,
      buf_acc_data_13_16_56_46_sva_mx0, buf_acc_data_13_17_56_46_sva_mx0, buf_acc_data_14_0_56_46_sva_mx0,
      buf_acc_data_14_1_56_46_sva_mx0, buf_acc_data_14_2_56_46_sva_mx0, buf_acc_data_14_3_56_46_sva_mx0,
      buf_acc_data_14_4_56_46_sva_mx0, buf_acc_data_14_5_56_46_sva_mx0, buf_acc_data_14_6_56_46_sva_mx0,
      buf_acc_data_14_7_56_46_sva_mx0, buf_acc_data_14_8_56_46_sva_mx0, buf_acc_data_14_9_56_46_sva_mx0,
      buf_acc_data_14_10_56_46_sva_mx0, buf_acc_data_14_11_56_46_sva_mx0, buf_acc_data_14_12_56_46_sva_mx0,
      buf_acc_data_14_13_56_46_sva_mx0, buf_acc_data_14_14_56_46_sva_mx0, buf_acc_data_14_15_56_46_sva_mx0,
      buf_acc_data_14_16_56_46_sva_mx0, buf_acc_data_14_17_56_46_sva_mx0, buf_acc_data_15_0_56_46_sva_mx0,
      buf_acc_data_15_1_56_46_sva_mx0, buf_acc_data_15_2_56_46_sva_mx0, buf_acc_data_15_3_56_46_sva_mx0,
      buf_acc_data_15_4_56_46_sva_mx0, buf_acc_data_15_5_56_46_sva_mx0, buf_acc_data_15_6_56_46_sva_mx0,
      buf_acc_data_15_7_56_46_sva_mx0, buf_acc_data_15_8_56_46_sva_mx0, buf_acc_data_15_9_56_46_sva_mx0,
      buf_acc_data_15_10_56_46_sva_mx0, buf_acc_data_15_11_56_46_sva_mx0, buf_acc_data_15_12_56_46_sva_mx0,
      buf_acc_data_15_13_56_46_sva_mx0, buf_acc_data_15_14_56_46_sva_mx0, buf_acc_data_15_15_56_46_sva_mx0,
      buf_acc_data_15_16_56_46_sva_mx0, buf_acc_data_15_17_56_46_sva_mx0, buf_acc_data_16_0_56_46_sva_mx0,
      buf_acc_data_16_1_56_46_sva_mx0, buf_acc_data_16_2_56_46_sva_mx0, buf_acc_data_16_3_56_46_sva_mx0,
      buf_acc_data_16_4_56_46_sva_mx0, buf_acc_data_16_5_56_46_sva_mx0, buf_acc_data_16_6_56_46_sva_mx0,
      buf_acc_data_16_7_56_46_sva_mx0, buf_acc_data_16_8_56_46_sva_mx0, buf_acc_data_16_9_56_46_sva_mx0,
      buf_acc_data_16_10_56_46_sva_mx0, buf_acc_data_16_11_56_46_sva_mx0, buf_acc_data_16_12_56_46_sva_mx0,
      buf_acc_data_16_13_56_46_sva_mx0, buf_acc_data_16_14_56_46_sva_mx0, buf_acc_data_16_15_56_46_sva_mx0,
      buf_acc_data_16_16_56_46_sva_mx0, buf_acc_data_16_17_56_46_sva_mx0, buf_acc_data_17_0_56_46_sva_mx0,
      buf_acc_data_17_1_56_46_sva_mx0, buf_acc_data_17_2_56_46_sva_mx0, buf_acc_data_17_3_56_46_sva_mx0,
      buf_acc_data_17_4_56_46_sva_mx0, buf_acc_data_17_5_56_46_sva_mx0, buf_acc_data_17_6_56_46_sva_mx0,
      buf_acc_data_17_7_56_46_sva_mx0, buf_acc_data_17_8_56_46_sva_mx0, buf_acc_data_17_9_56_46_sva_mx0,
      buf_acc_data_17_10_56_46_sva_mx0, buf_acc_data_17_11_56_46_sva_mx0, buf_acc_data_17_12_56_46_sva_mx0,
      buf_acc_data_17_13_56_46_sva_mx0, buf_acc_data_17_14_56_46_sva_mx0, buf_acc_data_17_15_56_46_sva_mx0,
      buf_acc_data_17_16_56_46_sva_mx0, buf_acc_data_17_17_56_46_sva_mx0, {CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3
      , CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_1_0});
  assign exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0 = exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2
      | (~(lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2 & CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_and_1_tmp));
  assign CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6 = MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2,
      CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_and_1_tmp);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2283_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1_mx0w0,
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1, and_765_cse);
  assign exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1 = CONVOLUTION_LOOP_for_for_for_for_mux_2283_nl
      & exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1;
  assign or_1135_tmp = (STORE_LOOP_or_tmp_1 & (~ dma_read_ctrl_rsci_irdy_mxwt)) |
      STORE_LOOP_or_2_itm_1;
  assign nor_390_nl = ~(STORE_LOOP_and_15_itm_1 | or_1135_tmp);
  assign and_917_nl = STORE_LOOP_and_15_itm_1 & (~ or_1135_tmp);
  assign LOAD_LOOP_i_lpi_2_dfm_2_mx0w0 = MUX1HOT_v_16_3_2((signext_16_1(~ dma_read_ctrl_rsci_irdy_mxwt)),
      LOAD_LOOP_i_sva_1_1, LOAD_LOOP_i_lpi_2, {nor_390_nl , and_917_nl , or_1135_tmp});
  assign STORE_LOOP_and_4_cse = exit_PADDING_LOOP_for_lpi_2_dfm_4 & STORE_LOOP_equal_tmp_5;
  assign PADDING_LOOP_for_for_mux_2_nl = MUX_s_1_2_2(PADDING_LOOP_for_for_and_psp_mx1w0,
      PADDING_LOOP_for_for_and_psp, mux_tmp_356);
  assign or_1142_nl = (STORE_LOOP_and_4_cse & exit_PADDING_LOOP_lpi_2_dfm_mx0w0 &
      PADDING_LOOP_for_for_and_psp_mx1w0) | (PADDING_LOOP_for_for_mux_2_nl & (~ exit_PADDING_LOOP_for_lpi_2_dfm_4)
      & STORE_LOOP_equal_tmp_5);
  assign mux_557_nl = MUX_v_5_2_2(PADDING_LOOP_for_row_4_0_lpi_2, PADDING_LOOP_for_row_4_0_sva_2,
      or_1142_nl);
  assign nor_398_nl = ~((STORE_LOOP_and_4_cse & (~ exit_PADDING_LOOP_lpi_2_dfm_mx0w0))
      | STORE_LOOP_and_30_cse);
  assign PADDING_LOOP_for_row_4_0_lpi_2_dfm_5_mx0w0 = MUX_v_5_2_2(5'b00000, mux_557_nl,
      nor_398_nl);
  assign LOAD_LOOP_LOAD_LOOP_and_2_nl = lfst_exit_PADDING_LOOP_for_lpi_2 & (~ exit_LOAD_LOOP_lpi_2_dfm_1);
  assign STORE_LOOP_or_2327_nl = STORE_LOOP_or_tmp_mx0w0 | STORE_LOOP_equal_tmp_2_mx0w0
      | STORE_LOOP_equal_tmp_4 | STORE_LOOP_or_tmp_2;
  assign lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0 = MUX1HOT_s_1_3_2(lfst_exit_PADDING_LOOP_for_lpi_2,
      LOAD_LOOP_LOAD_LOOP_and_2_nl, (~ exit_PADDING_LOOP_for_lpi_2_dfm_4), {STORE_LOOP_or_2327_nl
      , STORE_LOOP_equal_tmp_6 , STORE_LOOP_equal_tmp_5});
  assign and_876_tmp = (~((~(exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0 & or_dcpl_65))
      & exit_PADDING_LOOP_for_for_lpi_2_dfm_1)) & STORE_LOOP_equal_tmp_5;
  assign STORE_LOOP_and_6_tmp = exit_PADDING_LOOP_for_for_lpi_2_dfm_1 & STORE_LOOP_equal_tmp_5;
  assign PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_1_nl = MUX_v_5_2_2(5'b00000,
      PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5, exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0);
  assign nor_391_nl = ~(STORE_LOOP_and_6_tmp | and_876_tmp);
  assign and_915_nl = STORE_LOOP_and_6_tmp & (~ and_876_tmp);
  assign PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4_mx0w0 = MUX1HOT_v_5_3_2(PADDING_LOOP_for_for_col_4_0_lpi_2,
      PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_1_nl, PADDING_LOOP_for_for_col_4_0_sva_2,
      {nor_391_nl , and_915_nl , and_876_tmp});
  assign PADDING_LOOP_PADDING_LOOP_and_2_nl = lfst_exit_CONVOLUTION_LOOP_for_lpi_2
      & (~ exit_PADDING_LOOP_lpi_2_dfm_3);
  assign STORE_LOOP_or_2323_nl = STORE_LOOP_or_tmp_mx0w0 | STORE_LOOP_equal_tmp_6
      | STORE_LOOP_equal_tmp_4 | STORE_LOOP_or_tmp_2;
  assign lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0 = MUX1HOT_s_1_3_2(lfst_exit_CONVOLUTION_LOOP_for_lpi_2,
      PADDING_LOOP_PADDING_LOOP_and_2_nl, (~ exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4),
      {STORE_LOOP_or_2323_nl , STORE_LOOP_equal_tmp_5 , STORE_LOOP_equal_tmp_2_mx0w0});
  assign STORE_LOOP_and_9_m1c = (~ exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4) & STORE_LOOP_equal_tmp_2_mx0w0;
  assign STORE_LOOP_and_10_cse = exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4 & STORE_LOOP_equal_tmp_2_mx0w0;
  assign nor_384_m1c = ~(or_dcpl_162 | or_dcpl_163);
  assign and_907_nl = (~ STORE_LOOP_and_10_cse) & nor_384_m1c;
  assign and_908_nl = STORE_LOOP_and_10_cse & nor_384_m1c;
  assign CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5_mx0w0 = MUX1HOT_v_5_4_2(CONVOLUTION_LOOP_for_for_i_4_0_lpi_2,
      ({{4{exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0}}, exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0}),
      CONVOLUTION_LOOP_for_for_i_4_0_sva_2, CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6,
      {and_907_nl , and_908_nl , or_dcpl_162 , or_dcpl_163});
  assign STORE_LOOP_and_11_m1c = (~ exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3)
      & STORE_LOOP_equal_tmp_2_mx0w0;
  assign STORE_LOOP_and_12_cse = exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3 &
      STORE_LOOP_equal_tmp_2_mx0w0;
  assign nor_385_m1c = ~(or_dcpl_168 | or_dcpl_169);
  assign and_905_nl = (~ STORE_LOOP_and_12_cse) & nor_385_m1c;
  assign and_906_nl = STORE_LOOP_and_12_cse & nor_385_m1c;
  assign CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5_mx0w0 = MUX1HOT_v_5_4_2(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2,
      ({{4{exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0}}, exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0}),
      CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2, CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6,
      {and_905_nl , and_906_nl , or_dcpl_168 , or_dcpl_169});
  assign STORE_LOOP_nand_nl = ~(STORE_LOOP_equal_tmp_2_mx0w0 & (~((~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0)
      & STORE_LOOP_and_1_m1c_1)));
  assign STORE_LOOP_and_18_nl = exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0
      & STORE_LOOP_and_1_m1c_1;
  assign CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2_mx0w0 = MUX1HOT_v_8_3_2(CONVOLUTION_LOOP_for_for_for_x_lpi_2,
      (z_out_11_16_0[7:0]), z_out_13, {STORE_LOOP_nand_nl , STORE_LOOP_and_18_nl
      , STORE_LOOP_asn_3330});
  assign STORE_LOOP_and_25_nl = (~ CONVOLUTION_LOOP_for_for_for_for_for_and_5_tmp_1)
      & STORE_LOOP_equal_tmp_2_mx0w0;
  assign STORE_LOOP_and_26_nl = CONVOLUTION_LOOP_for_for_for_for_for_and_5_tmp_1
      & STORE_LOOP_equal_tmp_2_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3_mx0w0 = MUX1HOT_v_3_3_2(CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2,
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_4, CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2,
      {(~ STORE_LOOP_equal_tmp_2_mx0w0) , STORE_LOOP_and_25_nl , STORE_LOOP_and_26_nl});
  assign or_1156_tmp = (exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1_mx0w0 &
      or_1062_cse & STORE_LOOP_asn_3330) | STORE_LOOP_and_1_m1c_1;
  assign CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_and_nl
      = MUX_v_3_2_2(3'b000, CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_5,
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1_mx0w0);
  assign nor_392_nl = ~(STORE_LOOP_asn_3330 | or_1156_tmp);
  assign and_913_nl = STORE_LOOP_asn_3330 & (~ or_1156_tmp);
  assign CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4_mx0w0 = MUX1HOT_v_3_3_2(CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2,
      CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_and_nl,
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2, {nor_392_nl , and_913_nl
      , or_1156_tmp});
  assign or_1160_tmp = or_dcpl_135 | (exit_STORE_LOOP_sva_3 & STORE_LOOP_equal_tmp_4)
      | STORE_LOOP_and_33_cse | STORE_LOOP_equal_tmp_5 | STORE_LOOP_equal_tmp_6;
  assign STORE_LOOP_and_27_tmp = (~ exit_STORE_LOOP_sva_3) & STORE_LOOP_equal_tmp_4;
  assign nor_393_nl = ~(STORE_LOOP_and_27_tmp | or_1160_tmp);
  assign STORE_LOOP_i_13_0_lpi_2_dfm_2_mx0w0 = MUX1HOT_v_14_3_2((signext_14_1(~ exit_CONVOLUTION_LOOP_lpi_2_dfm_2_mx0w0)),
      STORE_LOOP_i_13_0_sva_2, STORE_LOOP_i_13_0_lpi_2, {nor_393_nl , STORE_LOOP_and_27_tmp
      , or_1160_tmp});
  assign STORE_LOOP_mux_31_nl = MUX_s_1_2_2(reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse,
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_5_1_2_cse, STORE_LOOP_and_35_itm_1);
  assign STORE_LOOP_STORE_LOOP_or_tmp = (STORE_LOOP_mux_31_nl & (~(STORE_LOOP_or_tmp_1
      | STORE_LOOP_and_30_itm_1))) | STORE_LOOP_and_32_itm_1 | STORE_LOOP_and_34_ssc_1;
  assign STORE_LOOP_mux1h_2331_nl = MUX1HOT_s_1_3_2((~ dma_read_ctrl_rsci_irdy_mxwt),
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse, reg_lfst_exit_STORE_LOOP_lpi_2_dfm_5_1_2_cse,
      {STORE_LOOP_or_tmp_1 , STORE_LOOP_or_2332_itm_1 , STORE_LOOP_and_35_itm_1});
  assign STORE_LOOP_or_2336_tmp = (STORE_LOOP_mux1h_2331_nl & (~ STORE_LOOP_and_32_itm_1))
      | STORE_LOOP_and_30_itm_1 | STORE_LOOP_and_34_ssc_1;
  assign STORE_LOOP_mux_34_nl = MUX_s_1_2_2(dma_read_ctrl_rsci_irdy_mxwt, reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse,
      STORE_LOOP_or_2332_itm_1);
  assign STORE_LOOP_or_2335_tmp = (STORE_LOOP_mux_34_nl & (~ STORE_LOOP_and_35_itm_1)
      & (~(STORE_LOOP_and_32_itm_1 | STORE_LOOP_and_34_ssc_1))) | STORE_LOOP_and_30_itm_1;
  assign nl_if_acc_4_cse_1 = ({(z_out_5_12_0[6:0]) , 1'b0}) - (conf_info_rsci_idat_mxwt[103:96]);
  assign if_acc_4_cse_1 = nl_if_acc_4_cse_1[7:0];
  assign nl_else_acc_2_psp_sva_1 = conv_u2s_10_11(z_out_2) + conv_s2s_9_11({1'b1
      , (conf_info_rsci_idat_mxwt[167:160])});
  assign else_acc_2_psp_sva_1 = nl_else_acc_2_psp_sva_1[10:0];
  assign nl_else_acc_psp_sva_1 = conv_u2s_10_11(z_out_2) + conv_s2s_9_11({1'b1 ,
      (conf_info_rsci_idat_mxwt[199:192])});
  assign else_acc_psp_sva_1 = nl_else_acc_psp_sva_1[10:0];
  assign LOAD_LOOP_i_lpi_2_mx1 = MUX_v_16_2_2(LOAD_LOOP_i_lpi_2_dfm_2_mx0w0, LOAD_LOOP_i_lpi_2,
      or_214_cse);
  assign CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1 = MUX_v_5_2_2(CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0,
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0, or_214_cse);
  assign nl_asn_3_mx0w1 = if_acc_4_cse_1 + (conf_info_rsci_idat_mxwt[199:192]) +
      8'b00000001;
  assign asn_3_mx0w1 = nl_asn_3_mx0w1[7:0];
  assign operator_42_true_1_and_nl = (else_acc_2_psp_sva_1[10]) & (else_acc_2_psp_sva_1[0]);
  assign nl_asn_1_mx0w0 = (else_acc_2_psp_sva_1[8:1]) + conv_u2u_1_8(operator_42_true_1_and_nl)
      + 8'b00000001;
  assign asn_1_mx0w0 = nl_asn_1_mx0w0[7:0];
  assign nl_asn_mx0w1 = if_acc_4_cse_1 + (conf_info_rsci_idat_mxwt[167:160]) + 8'b00000001;
  assign asn_mx0w1 = nl_asn_mx0w1[7:0];
  assign STORE_LOOP_STORE_LOOP_nor_2_nl = ~(STORE_LOOP_STORE_LOOP_or_tmp | STORE_LOOP_or_2335_tmp
      | STORE_LOOP_or_2336_tmp);
  assign or_789_nl = BATCH_LOOP_asn_itm_1 | exit_BATCH_LOOP_lpi_2_dfm_2_1 | (~ BATCH_LOOP_and_4_tmp);
  assign exitL_exit_STORE_LOOP_sva_mx1 = MUX_s_1_2_2(STORE_LOOP_STORE_LOOP_nor_2_nl,
      exitL_exit_STORE_LOOP_sva, or_789_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2296_nl = MUX_s_1_2_2(buf_acc_data_17_17_0_sva,
      buf_acc_data_17_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2296_nl,
      buf_acc_data_17_17_0_sva, or_dcpl_124);
  assign buf_acc_data_17_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_17_45_1_sva_dfm_1,
      buf_acc_data_17_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_17_56_46_sva_dfm_1,
      buf_acc_data_17_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2298_nl = MUX_s_1_2_2(buf_acc_data_0_0_0_sva,
      buf_acc_data_0_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2298_nl,
      buf_acc_data_0_0_0_sva, or_dcpl_124);
  assign buf_acc_data_0_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_0_45_1_sva_dfm_1,
      buf_acc_data_0_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_0_56_46_sva_dfm_1,
      buf_acc_data_0_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2300_nl = MUX_s_1_2_2(buf_acc_data_17_16_0_sva,
      buf_acc_data_17_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2300_nl,
      buf_acc_data_17_16_0_sva, or_dcpl_124);
  assign buf_acc_data_17_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_16_45_1_sva_dfm_1,
      buf_acc_data_17_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_16_56_46_sva_dfm_1,
      buf_acc_data_17_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2302_nl = MUX_s_1_2_2(buf_acc_data_0_1_0_sva,
      buf_acc_data_0_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2302_nl,
      buf_acc_data_0_1_0_sva, or_dcpl_124);
  assign buf_acc_data_0_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_1_45_1_sva_dfm_1,
      buf_acc_data_0_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_1_56_46_sva_dfm_1,
      buf_acc_data_0_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2304_nl = MUX_s_1_2_2(buf_acc_data_17_15_0_sva,
      buf_acc_data_17_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2304_nl,
      buf_acc_data_17_15_0_sva, or_dcpl_124);
  assign buf_acc_data_17_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_15_45_1_sva_dfm_1,
      buf_acc_data_17_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_15_56_46_sva_dfm_1,
      buf_acc_data_17_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2306_nl = MUX_s_1_2_2(buf_acc_data_0_2_0_sva,
      buf_acc_data_0_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2306_nl,
      buf_acc_data_0_2_0_sva, or_dcpl_124);
  assign buf_acc_data_0_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_2_45_1_sva_dfm_1,
      buf_acc_data_0_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_2_56_46_sva_dfm_1,
      buf_acc_data_0_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2308_nl = MUX_s_1_2_2(buf_acc_data_17_14_0_sva,
      buf_acc_data_17_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2308_nl,
      buf_acc_data_17_14_0_sva, or_dcpl_124);
  assign buf_acc_data_17_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_14_45_1_sva_dfm_1,
      buf_acc_data_17_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_14_56_46_sva_dfm_1,
      buf_acc_data_17_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2310_nl = MUX_s_1_2_2(buf_acc_data_0_3_0_sva,
      buf_acc_data_0_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2310_nl,
      buf_acc_data_0_3_0_sva, or_dcpl_124);
  assign buf_acc_data_0_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_3_45_1_sva_dfm_1,
      buf_acc_data_0_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_3_56_46_sva_dfm_1,
      buf_acc_data_0_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2312_nl = MUX_s_1_2_2(buf_acc_data_17_13_0_sva,
      buf_acc_data_17_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2312_nl,
      buf_acc_data_17_13_0_sva, or_dcpl_124);
  assign buf_acc_data_17_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_13_45_1_sva_dfm_1,
      buf_acc_data_17_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_13_56_46_sva_dfm_1,
      buf_acc_data_17_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2314_nl = MUX_s_1_2_2(buf_acc_data_0_4_0_sva,
      buf_acc_data_0_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2314_nl,
      buf_acc_data_0_4_0_sva, or_dcpl_124);
  assign buf_acc_data_0_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_4_45_1_sva_dfm_1,
      buf_acc_data_0_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_4_56_46_sva_dfm_1,
      buf_acc_data_0_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2316_nl = MUX_s_1_2_2(buf_acc_data_17_12_0_sva,
      buf_acc_data_17_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2316_nl,
      buf_acc_data_17_12_0_sva, or_dcpl_124);
  assign buf_acc_data_17_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_12_45_1_sva_dfm_1,
      buf_acc_data_17_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_12_56_46_sva_dfm_1,
      buf_acc_data_17_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2318_nl = MUX_s_1_2_2(buf_acc_data_0_5_0_sva,
      buf_acc_data_0_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2318_nl,
      buf_acc_data_0_5_0_sva, or_dcpl_124);
  assign buf_acc_data_0_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_5_45_1_sva_dfm_1,
      buf_acc_data_0_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_5_56_46_sva_dfm_1,
      buf_acc_data_0_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2320_nl = MUX_s_1_2_2(buf_acc_data_17_11_0_sva,
      buf_acc_data_17_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2320_nl,
      buf_acc_data_17_11_0_sva, or_dcpl_124);
  assign buf_acc_data_17_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_11_45_1_sva_dfm_1,
      buf_acc_data_17_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_11_56_46_sva_dfm_1,
      buf_acc_data_17_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2322_nl = MUX_s_1_2_2(buf_acc_data_0_6_0_sva,
      buf_acc_data_0_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2322_nl,
      buf_acc_data_0_6_0_sva, or_dcpl_124);
  assign buf_acc_data_0_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_6_45_1_sva_dfm_1,
      buf_acc_data_0_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_6_56_46_sva_dfm_1,
      buf_acc_data_0_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2324_nl = MUX_s_1_2_2(buf_acc_data_17_10_0_sva,
      buf_acc_data_17_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2324_nl,
      buf_acc_data_17_10_0_sva, or_dcpl_124);
  assign buf_acc_data_17_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_10_45_1_sva_dfm_1,
      buf_acc_data_17_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_10_56_46_sva_dfm_1,
      buf_acc_data_17_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2326_nl = MUX_s_1_2_2(buf_acc_data_0_7_0_sva,
      buf_acc_data_0_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2326_nl,
      buf_acc_data_0_7_0_sva, or_dcpl_124);
  assign buf_acc_data_0_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_7_45_1_sva_dfm_1,
      buf_acc_data_0_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_7_56_46_sva_dfm_1,
      buf_acc_data_0_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2328_nl = MUX_s_1_2_2(buf_acc_data_17_9_0_sva,
      buf_acc_data_17_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2328_nl,
      buf_acc_data_17_9_0_sva, or_dcpl_124);
  assign buf_acc_data_17_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_9_45_1_sva_dfm_1,
      buf_acc_data_17_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_9_56_46_sva_dfm_1,
      buf_acc_data_17_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2330_nl = MUX_s_1_2_2(buf_acc_data_0_8_0_sva,
      buf_acc_data_0_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2330_nl,
      buf_acc_data_0_8_0_sva, or_dcpl_124);
  assign buf_acc_data_0_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_8_45_1_sva_dfm_1,
      buf_acc_data_0_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_8_56_46_sva_dfm_1,
      buf_acc_data_0_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2332_nl = MUX_s_1_2_2(buf_acc_data_17_8_0_sva,
      buf_acc_data_17_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2332_nl,
      buf_acc_data_17_8_0_sva, or_dcpl_124);
  assign buf_acc_data_17_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_8_45_1_sva_dfm_1,
      buf_acc_data_17_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_8_56_46_sva_dfm_1,
      buf_acc_data_17_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2334_nl = MUX_s_1_2_2(buf_acc_data_0_9_0_sva,
      buf_acc_data_0_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2334_nl,
      buf_acc_data_0_9_0_sva, or_dcpl_124);
  assign buf_acc_data_0_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_9_45_1_sva_dfm_1,
      buf_acc_data_0_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_9_56_46_sva_dfm_1,
      buf_acc_data_0_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2336_nl = MUX_s_1_2_2(buf_acc_data_17_7_0_sva,
      buf_acc_data_17_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2336_nl,
      buf_acc_data_17_7_0_sva, or_dcpl_124);
  assign buf_acc_data_17_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_7_45_1_sva_dfm_1,
      buf_acc_data_17_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_7_56_46_sva_dfm_1,
      buf_acc_data_17_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2338_nl = MUX_s_1_2_2(buf_acc_data_0_10_0_sva,
      buf_acc_data_0_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2338_nl,
      buf_acc_data_0_10_0_sva, or_dcpl_124);
  assign buf_acc_data_0_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_10_45_1_sva_dfm_1,
      buf_acc_data_0_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_10_56_46_sva_dfm_1,
      buf_acc_data_0_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2340_nl = MUX_s_1_2_2(buf_acc_data_17_6_0_sva,
      buf_acc_data_17_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2340_nl,
      buf_acc_data_17_6_0_sva, or_dcpl_124);
  assign buf_acc_data_17_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_6_45_1_sva_dfm_1,
      buf_acc_data_17_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_6_56_46_sva_dfm_1,
      buf_acc_data_17_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2342_nl = MUX_s_1_2_2(buf_acc_data_0_11_0_sva,
      buf_acc_data_0_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2342_nl,
      buf_acc_data_0_11_0_sva, or_dcpl_124);
  assign buf_acc_data_0_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_11_45_1_sva_dfm_1,
      buf_acc_data_0_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_11_56_46_sva_dfm_1,
      buf_acc_data_0_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2344_nl = MUX_s_1_2_2(buf_acc_data_17_5_0_sva,
      buf_acc_data_17_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2344_nl,
      buf_acc_data_17_5_0_sva, or_dcpl_124);
  assign buf_acc_data_17_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_5_45_1_sva_dfm_1,
      buf_acc_data_17_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_5_56_46_sva_dfm_1,
      buf_acc_data_17_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2346_nl = MUX_s_1_2_2(buf_acc_data_0_12_0_sva,
      buf_acc_data_0_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2346_nl,
      buf_acc_data_0_12_0_sva, or_dcpl_124);
  assign buf_acc_data_0_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_12_45_1_sva_dfm_1,
      buf_acc_data_0_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_12_56_46_sva_dfm_1,
      buf_acc_data_0_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2348_nl = MUX_s_1_2_2(buf_acc_data_17_4_0_sva,
      buf_acc_data_17_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2348_nl,
      buf_acc_data_17_4_0_sva, or_dcpl_124);
  assign buf_acc_data_17_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_4_45_1_sva_dfm_1,
      buf_acc_data_17_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_4_56_46_sva_dfm_1,
      buf_acc_data_17_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2350_nl = MUX_s_1_2_2(buf_acc_data_0_13_0_sva,
      buf_acc_data_0_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2350_nl,
      buf_acc_data_0_13_0_sva, or_dcpl_124);
  assign buf_acc_data_0_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_13_45_1_sva_dfm_1,
      buf_acc_data_0_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_13_56_46_sva_dfm_1,
      buf_acc_data_0_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2352_nl = MUX_s_1_2_2(buf_acc_data_17_3_0_sva,
      buf_acc_data_17_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2352_nl,
      buf_acc_data_17_3_0_sva, or_dcpl_124);
  assign buf_acc_data_17_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_3_45_1_sva_dfm_1,
      buf_acc_data_17_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_3_56_46_sva_dfm_1,
      buf_acc_data_17_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2354_nl = MUX_s_1_2_2(buf_acc_data_0_14_0_sva,
      buf_acc_data_0_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2354_nl,
      buf_acc_data_0_14_0_sva, or_dcpl_124);
  assign buf_acc_data_0_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_14_45_1_sva_dfm_1,
      buf_acc_data_0_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_14_56_46_sva_dfm_1,
      buf_acc_data_0_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2356_nl = MUX_s_1_2_2(buf_acc_data_17_2_0_sva,
      buf_acc_data_17_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2356_nl,
      buf_acc_data_17_2_0_sva, or_dcpl_124);
  assign buf_acc_data_17_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_2_45_1_sva_dfm_1,
      buf_acc_data_17_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_2_56_46_sva_dfm_1,
      buf_acc_data_17_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2358_nl = MUX_s_1_2_2(buf_acc_data_0_15_0_sva,
      buf_acc_data_0_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2358_nl,
      buf_acc_data_0_15_0_sva, or_dcpl_124);
  assign buf_acc_data_0_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_15_45_1_sva_dfm_1,
      buf_acc_data_0_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_15_56_46_sva_dfm_1,
      buf_acc_data_0_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2360_nl = MUX_s_1_2_2(buf_acc_data_17_1_0_sva,
      buf_acc_data_17_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2360_nl,
      buf_acc_data_17_1_0_sva, or_dcpl_124);
  assign buf_acc_data_17_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_1_45_1_sva_dfm_1,
      buf_acc_data_17_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_1_56_46_sva_dfm_1,
      buf_acc_data_17_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2362_nl = MUX_s_1_2_2(buf_acc_data_0_16_0_sva,
      buf_acc_data_0_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2362_nl,
      buf_acc_data_0_16_0_sva, or_dcpl_124);
  assign buf_acc_data_0_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_16_45_1_sva_dfm_1,
      buf_acc_data_0_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_16_56_46_sva_dfm_1,
      buf_acc_data_0_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2364_nl = MUX_s_1_2_2(buf_acc_data_17_0_0_sva,
      buf_acc_data_17_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_17_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2364_nl,
      buf_acc_data_17_0_0_sva, or_dcpl_124);
  assign buf_acc_data_17_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_17_0_45_1_sva_dfm_1,
      buf_acc_data_17_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_17_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_17_0_56_46_sva_dfm_1,
      buf_acc_data_17_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2366_nl = MUX_s_1_2_2(buf_acc_data_0_17_0_sva,
      buf_acc_data_0_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_0_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2366_nl,
      buf_acc_data_0_17_0_sva, or_dcpl_124);
  assign buf_acc_data_0_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_0_17_45_1_sva_dfm_1,
      buf_acc_data_0_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_0_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_0_17_56_46_sva_dfm_1,
      buf_acc_data_0_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2368_nl = MUX_s_1_2_2(buf_acc_data_16_17_0_sva,
      buf_acc_data_16_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2368_nl,
      buf_acc_data_16_17_0_sva, or_dcpl_124);
  assign buf_acc_data_16_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_17_45_1_sva_dfm_1,
      buf_acc_data_16_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_17_56_46_sva_dfm_1,
      buf_acc_data_16_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2370_nl = MUX_s_1_2_2(buf_acc_data_1_0_0_sva,
      buf_acc_data_1_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2370_nl,
      buf_acc_data_1_0_0_sva, or_dcpl_124);
  assign buf_acc_data_1_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_0_45_1_sva_dfm_1,
      buf_acc_data_1_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_0_56_46_sva_dfm_1,
      buf_acc_data_1_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2372_nl = MUX_s_1_2_2(buf_acc_data_16_16_0_sva,
      buf_acc_data_16_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2372_nl,
      buf_acc_data_16_16_0_sva, or_dcpl_124);
  assign buf_acc_data_16_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_16_45_1_sva_dfm_1,
      buf_acc_data_16_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_16_56_46_sva_dfm_1,
      buf_acc_data_16_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2374_nl = MUX_s_1_2_2(buf_acc_data_1_1_0_sva,
      buf_acc_data_1_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2374_nl,
      buf_acc_data_1_1_0_sva, or_dcpl_124);
  assign buf_acc_data_1_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_1_45_1_sva_dfm_1,
      buf_acc_data_1_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_1_56_46_sva_dfm_1,
      buf_acc_data_1_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2376_nl = MUX_s_1_2_2(buf_acc_data_16_15_0_sva,
      buf_acc_data_16_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2376_nl,
      buf_acc_data_16_15_0_sva, or_dcpl_124);
  assign buf_acc_data_16_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_15_45_1_sva_dfm_1,
      buf_acc_data_16_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_15_56_46_sva_dfm_1,
      buf_acc_data_16_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2378_nl = MUX_s_1_2_2(buf_acc_data_1_2_0_sva,
      buf_acc_data_1_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2378_nl,
      buf_acc_data_1_2_0_sva, or_dcpl_124);
  assign buf_acc_data_1_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_2_45_1_sva_dfm_1,
      buf_acc_data_1_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_2_56_46_sva_dfm_1,
      buf_acc_data_1_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2380_nl = MUX_s_1_2_2(buf_acc_data_16_14_0_sva,
      buf_acc_data_16_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2380_nl,
      buf_acc_data_16_14_0_sva, or_dcpl_124);
  assign buf_acc_data_16_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_14_45_1_sva_dfm_1,
      buf_acc_data_16_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_14_56_46_sva_dfm_1,
      buf_acc_data_16_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2382_nl = MUX_s_1_2_2(buf_acc_data_1_3_0_sva,
      buf_acc_data_1_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2382_nl,
      buf_acc_data_1_3_0_sva, or_dcpl_124);
  assign buf_acc_data_1_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_3_45_1_sva_dfm_1,
      buf_acc_data_1_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_3_56_46_sva_dfm_1,
      buf_acc_data_1_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2384_nl = MUX_s_1_2_2(buf_acc_data_16_13_0_sva,
      buf_acc_data_16_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2384_nl,
      buf_acc_data_16_13_0_sva, or_dcpl_124);
  assign buf_acc_data_16_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_13_45_1_sva_dfm_1,
      buf_acc_data_16_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_13_56_46_sva_dfm_1,
      buf_acc_data_16_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2386_nl = MUX_s_1_2_2(buf_acc_data_1_4_0_sva,
      buf_acc_data_1_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2386_nl,
      buf_acc_data_1_4_0_sva, or_dcpl_124);
  assign buf_acc_data_1_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_4_45_1_sva_dfm_1,
      buf_acc_data_1_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_4_56_46_sva_dfm_1,
      buf_acc_data_1_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2388_nl = MUX_s_1_2_2(buf_acc_data_16_12_0_sva,
      buf_acc_data_16_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2388_nl,
      buf_acc_data_16_12_0_sva, or_dcpl_124);
  assign buf_acc_data_16_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_12_45_1_sva_dfm_1,
      buf_acc_data_16_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_12_56_46_sva_dfm_1,
      buf_acc_data_16_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2390_nl = MUX_s_1_2_2(buf_acc_data_1_5_0_sva,
      buf_acc_data_1_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2390_nl,
      buf_acc_data_1_5_0_sva, or_dcpl_124);
  assign buf_acc_data_1_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_5_45_1_sva_dfm_1,
      buf_acc_data_1_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_5_56_46_sva_dfm_1,
      buf_acc_data_1_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2392_nl = MUX_s_1_2_2(buf_acc_data_16_11_0_sva,
      buf_acc_data_16_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2392_nl,
      buf_acc_data_16_11_0_sva, or_dcpl_124);
  assign buf_acc_data_16_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_11_45_1_sva_dfm_1,
      buf_acc_data_16_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_11_56_46_sva_dfm_1,
      buf_acc_data_16_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2394_nl = MUX_s_1_2_2(buf_acc_data_1_6_0_sva,
      buf_acc_data_1_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2394_nl,
      buf_acc_data_1_6_0_sva, or_dcpl_124);
  assign buf_acc_data_1_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_6_45_1_sva_dfm_1,
      buf_acc_data_1_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_6_56_46_sva_dfm_1,
      buf_acc_data_1_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2396_nl = MUX_s_1_2_2(buf_acc_data_16_10_0_sva,
      buf_acc_data_16_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2396_nl,
      buf_acc_data_16_10_0_sva, or_dcpl_124);
  assign buf_acc_data_16_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_10_45_1_sva_dfm_1,
      buf_acc_data_16_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_10_56_46_sva_dfm_1,
      buf_acc_data_16_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2398_nl = MUX_s_1_2_2(buf_acc_data_1_7_0_sva,
      buf_acc_data_1_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2398_nl,
      buf_acc_data_1_7_0_sva, or_dcpl_124);
  assign buf_acc_data_1_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_7_45_1_sva_dfm_1,
      buf_acc_data_1_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_7_56_46_sva_dfm_1,
      buf_acc_data_1_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2400_nl = MUX_s_1_2_2(buf_acc_data_16_9_0_sva,
      buf_acc_data_16_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2400_nl,
      buf_acc_data_16_9_0_sva, or_dcpl_124);
  assign buf_acc_data_16_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_9_45_1_sva_dfm_1,
      buf_acc_data_16_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_9_56_46_sva_dfm_1,
      buf_acc_data_16_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2402_nl = MUX_s_1_2_2(buf_acc_data_1_8_0_sva,
      buf_acc_data_1_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2402_nl,
      buf_acc_data_1_8_0_sva, or_dcpl_124);
  assign buf_acc_data_1_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_8_45_1_sva_dfm_1,
      buf_acc_data_1_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_8_56_46_sva_dfm_1,
      buf_acc_data_1_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2404_nl = MUX_s_1_2_2(buf_acc_data_16_8_0_sva,
      buf_acc_data_16_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2404_nl,
      buf_acc_data_16_8_0_sva, or_dcpl_124);
  assign buf_acc_data_16_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_8_45_1_sva_dfm_1,
      buf_acc_data_16_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_8_56_46_sva_dfm_1,
      buf_acc_data_16_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2406_nl = MUX_s_1_2_2(buf_acc_data_1_9_0_sva,
      buf_acc_data_1_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2406_nl,
      buf_acc_data_1_9_0_sva, or_dcpl_124);
  assign buf_acc_data_1_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_9_45_1_sva_dfm_1,
      buf_acc_data_1_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_9_56_46_sva_dfm_1,
      buf_acc_data_1_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2408_nl = MUX_s_1_2_2(buf_acc_data_16_7_0_sva,
      buf_acc_data_16_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2408_nl,
      buf_acc_data_16_7_0_sva, or_dcpl_124);
  assign buf_acc_data_16_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_7_45_1_sva_dfm_1,
      buf_acc_data_16_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_7_56_46_sva_dfm_1,
      buf_acc_data_16_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2410_nl = MUX_s_1_2_2(buf_acc_data_1_10_0_sva,
      buf_acc_data_1_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2410_nl,
      buf_acc_data_1_10_0_sva, or_dcpl_124);
  assign buf_acc_data_1_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_10_45_1_sva_dfm_1,
      buf_acc_data_1_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_10_56_46_sva_dfm_1,
      buf_acc_data_1_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2412_nl = MUX_s_1_2_2(buf_acc_data_16_6_0_sva,
      buf_acc_data_16_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2412_nl,
      buf_acc_data_16_6_0_sva, or_dcpl_124);
  assign buf_acc_data_16_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_6_45_1_sva_dfm_1,
      buf_acc_data_16_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_6_56_46_sva_dfm_1,
      buf_acc_data_16_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2414_nl = MUX_s_1_2_2(buf_acc_data_1_11_0_sva,
      buf_acc_data_1_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2414_nl,
      buf_acc_data_1_11_0_sva, or_dcpl_124);
  assign buf_acc_data_1_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_11_45_1_sva_dfm_1,
      buf_acc_data_1_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_11_56_46_sva_dfm_1,
      buf_acc_data_1_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2416_nl = MUX_s_1_2_2(buf_acc_data_16_5_0_sva,
      buf_acc_data_16_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2416_nl,
      buf_acc_data_16_5_0_sva, or_dcpl_124);
  assign buf_acc_data_16_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_5_45_1_sva_dfm_1,
      buf_acc_data_16_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_5_56_46_sva_dfm_1,
      buf_acc_data_16_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2418_nl = MUX_s_1_2_2(buf_acc_data_1_12_0_sva,
      buf_acc_data_1_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2418_nl,
      buf_acc_data_1_12_0_sva, or_dcpl_124);
  assign buf_acc_data_1_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_12_45_1_sva_dfm_1,
      buf_acc_data_1_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_12_56_46_sva_dfm_1,
      buf_acc_data_1_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2420_nl = MUX_s_1_2_2(buf_acc_data_16_4_0_sva,
      buf_acc_data_16_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2420_nl,
      buf_acc_data_16_4_0_sva, or_dcpl_124);
  assign buf_acc_data_16_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_4_45_1_sva_dfm_1,
      buf_acc_data_16_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_4_56_46_sva_dfm_1,
      buf_acc_data_16_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2422_nl = MUX_s_1_2_2(buf_acc_data_1_13_0_sva,
      buf_acc_data_1_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2422_nl,
      buf_acc_data_1_13_0_sva, or_dcpl_124);
  assign buf_acc_data_1_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_13_45_1_sva_dfm_1,
      buf_acc_data_1_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_13_56_46_sva_dfm_1,
      buf_acc_data_1_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2424_nl = MUX_s_1_2_2(buf_acc_data_16_3_0_sva,
      buf_acc_data_16_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2424_nl,
      buf_acc_data_16_3_0_sva, or_dcpl_124);
  assign buf_acc_data_16_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_3_45_1_sva_dfm_1,
      buf_acc_data_16_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_3_56_46_sva_dfm_1,
      buf_acc_data_16_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2426_nl = MUX_s_1_2_2(buf_acc_data_1_14_0_sva,
      buf_acc_data_1_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2426_nl,
      buf_acc_data_1_14_0_sva, or_dcpl_124);
  assign buf_acc_data_1_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_14_45_1_sva_dfm_1,
      buf_acc_data_1_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_14_56_46_sva_dfm_1,
      buf_acc_data_1_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2428_nl = MUX_s_1_2_2(buf_acc_data_16_2_0_sva,
      buf_acc_data_16_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2428_nl,
      buf_acc_data_16_2_0_sva, or_dcpl_124);
  assign buf_acc_data_16_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_2_45_1_sva_dfm_1,
      buf_acc_data_16_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_2_56_46_sva_dfm_1,
      buf_acc_data_16_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2430_nl = MUX_s_1_2_2(buf_acc_data_1_15_0_sva,
      buf_acc_data_1_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2430_nl,
      buf_acc_data_1_15_0_sva, or_dcpl_124);
  assign buf_acc_data_1_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_15_45_1_sva_dfm_1,
      buf_acc_data_1_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_15_56_46_sva_dfm_1,
      buf_acc_data_1_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2432_nl = MUX_s_1_2_2(buf_acc_data_16_1_0_sva,
      buf_acc_data_16_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2432_nl,
      buf_acc_data_16_1_0_sva, or_dcpl_124);
  assign buf_acc_data_16_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_1_45_1_sva_dfm_1,
      buf_acc_data_16_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_1_56_46_sva_dfm_1,
      buf_acc_data_16_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2434_nl = MUX_s_1_2_2(buf_acc_data_1_16_0_sva,
      buf_acc_data_1_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2434_nl,
      buf_acc_data_1_16_0_sva, or_dcpl_124);
  assign buf_acc_data_1_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_16_45_1_sva_dfm_1,
      buf_acc_data_1_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_16_56_46_sva_dfm_1,
      buf_acc_data_1_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2436_nl = MUX_s_1_2_2(buf_acc_data_16_0_0_sva,
      buf_acc_data_16_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_16_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2436_nl,
      buf_acc_data_16_0_0_sva, or_dcpl_124);
  assign buf_acc_data_16_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_16_0_45_1_sva_dfm_1,
      buf_acc_data_16_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_16_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_16_0_56_46_sva_dfm_1,
      buf_acc_data_16_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2438_nl = MUX_s_1_2_2(buf_acc_data_1_17_0_sva,
      buf_acc_data_1_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_1_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2438_nl,
      buf_acc_data_1_17_0_sva, or_dcpl_124);
  assign buf_acc_data_1_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_1_17_45_1_sva_dfm_1,
      buf_acc_data_1_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_1_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_1_17_56_46_sva_dfm_1,
      buf_acc_data_1_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2440_nl = MUX_s_1_2_2(buf_acc_data_15_17_0_sva,
      buf_acc_data_15_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2440_nl,
      buf_acc_data_15_17_0_sva, or_dcpl_124);
  assign buf_acc_data_15_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_17_45_1_sva_dfm_1,
      buf_acc_data_15_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_17_56_46_sva_dfm_1,
      buf_acc_data_15_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2442_nl = MUX_s_1_2_2(buf_acc_data_2_0_0_sva,
      buf_acc_data_2_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2442_nl,
      buf_acc_data_2_0_0_sva, or_dcpl_124);
  assign buf_acc_data_2_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_0_45_1_sva_dfm_1,
      buf_acc_data_2_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_0_56_46_sva_dfm_1,
      buf_acc_data_2_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2444_nl = MUX_s_1_2_2(buf_acc_data_15_16_0_sva,
      buf_acc_data_15_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2444_nl,
      buf_acc_data_15_16_0_sva, or_dcpl_124);
  assign buf_acc_data_15_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_16_45_1_sva_dfm_1,
      buf_acc_data_15_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_16_56_46_sva_dfm_1,
      buf_acc_data_15_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2446_nl = MUX_s_1_2_2(buf_acc_data_2_1_0_sva,
      buf_acc_data_2_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2446_nl,
      buf_acc_data_2_1_0_sva, or_dcpl_124);
  assign buf_acc_data_2_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_1_45_1_sva_dfm_1,
      buf_acc_data_2_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_1_56_46_sva_dfm_1,
      buf_acc_data_2_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2448_nl = MUX_s_1_2_2(buf_acc_data_15_15_0_sva,
      buf_acc_data_15_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2448_nl,
      buf_acc_data_15_15_0_sva, or_dcpl_124);
  assign buf_acc_data_15_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_15_45_1_sva_dfm_1,
      buf_acc_data_15_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_15_56_46_sva_dfm_1,
      buf_acc_data_15_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2450_nl = MUX_s_1_2_2(buf_acc_data_2_2_0_sva,
      buf_acc_data_2_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2450_nl,
      buf_acc_data_2_2_0_sva, or_dcpl_124);
  assign buf_acc_data_2_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_2_45_1_sva_dfm_1,
      buf_acc_data_2_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_2_56_46_sva_dfm_1,
      buf_acc_data_2_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2452_nl = MUX_s_1_2_2(buf_acc_data_15_14_0_sva,
      buf_acc_data_15_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2452_nl,
      buf_acc_data_15_14_0_sva, or_dcpl_124);
  assign buf_acc_data_15_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_14_45_1_sva_dfm_1,
      buf_acc_data_15_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_14_56_46_sva_dfm_1,
      buf_acc_data_15_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2454_nl = MUX_s_1_2_2(buf_acc_data_2_3_0_sva,
      buf_acc_data_2_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2454_nl,
      buf_acc_data_2_3_0_sva, or_dcpl_124);
  assign buf_acc_data_2_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_3_45_1_sva_dfm_1,
      buf_acc_data_2_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_3_56_46_sva_dfm_1,
      buf_acc_data_2_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2456_nl = MUX_s_1_2_2(buf_acc_data_15_13_0_sva,
      buf_acc_data_15_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2456_nl,
      buf_acc_data_15_13_0_sva, or_dcpl_124);
  assign buf_acc_data_15_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_13_45_1_sva_dfm_1,
      buf_acc_data_15_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_13_56_46_sva_dfm_1,
      buf_acc_data_15_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2458_nl = MUX_s_1_2_2(buf_acc_data_2_4_0_sva,
      buf_acc_data_2_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2458_nl,
      buf_acc_data_2_4_0_sva, or_dcpl_124);
  assign buf_acc_data_2_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_4_45_1_sva_dfm_1,
      buf_acc_data_2_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_4_56_46_sva_dfm_1,
      buf_acc_data_2_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2460_nl = MUX_s_1_2_2(buf_acc_data_15_12_0_sva,
      buf_acc_data_15_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2460_nl,
      buf_acc_data_15_12_0_sva, or_dcpl_124);
  assign buf_acc_data_15_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_12_45_1_sva_dfm_1,
      buf_acc_data_15_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_12_56_46_sva_dfm_1,
      buf_acc_data_15_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2462_nl = MUX_s_1_2_2(buf_acc_data_2_5_0_sva,
      buf_acc_data_2_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2462_nl,
      buf_acc_data_2_5_0_sva, or_dcpl_124);
  assign buf_acc_data_2_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_5_45_1_sva_dfm_1,
      buf_acc_data_2_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_5_56_46_sva_dfm_1,
      buf_acc_data_2_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2464_nl = MUX_s_1_2_2(buf_acc_data_15_11_0_sva,
      buf_acc_data_15_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2464_nl,
      buf_acc_data_15_11_0_sva, or_dcpl_124);
  assign buf_acc_data_15_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_11_45_1_sva_dfm_1,
      buf_acc_data_15_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_11_56_46_sva_dfm_1,
      buf_acc_data_15_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2466_nl = MUX_s_1_2_2(buf_acc_data_2_6_0_sva,
      buf_acc_data_2_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2466_nl,
      buf_acc_data_2_6_0_sva, or_dcpl_124);
  assign buf_acc_data_2_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_6_45_1_sva_dfm_1,
      buf_acc_data_2_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_6_56_46_sva_dfm_1,
      buf_acc_data_2_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2468_nl = MUX_s_1_2_2(buf_acc_data_15_10_0_sva,
      buf_acc_data_15_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2468_nl,
      buf_acc_data_15_10_0_sva, or_dcpl_124);
  assign buf_acc_data_15_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_10_45_1_sva_dfm_1,
      buf_acc_data_15_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_10_56_46_sva_dfm_1,
      buf_acc_data_15_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2470_nl = MUX_s_1_2_2(buf_acc_data_2_7_0_sva,
      buf_acc_data_2_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2470_nl,
      buf_acc_data_2_7_0_sva, or_dcpl_124);
  assign buf_acc_data_2_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_7_45_1_sva_dfm_1,
      buf_acc_data_2_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_7_56_46_sva_dfm_1,
      buf_acc_data_2_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2472_nl = MUX_s_1_2_2(buf_acc_data_15_9_0_sva,
      buf_acc_data_15_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2472_nl,
      buf_acc_data_15_9_0_sva, or_dcpl_124);
  assign buf_acc_data_15_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_9_45_1_sva_dfm_1,
      buf_acc_data_15_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_9_56_46_sva_dfm_1,
      buf_acc_data_15_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2474_nl = MUX_s_1_2_2(buf_acc_data_2_8_0_sva,
      buf_acc_data_2_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2474_nl,
      buf_acc_data_2_8_0_sva, or_dcpl_124);
  assign buf_acc_data_2_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_8_45_1_sva_dfm_1,
      buf_acc_data_2_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_8_56_46_sva_dfm_1,
      buf_acc_data_2_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2476_nl = MUX_s_1_2_2(buf_acc_data_15_8_0_sva,
      buf_acc_data_15_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2476_nl,
      buf_acc_data_15_8_0_sva, or_dcpl_124);
  assign buf_acc_data_15_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_8_45_1_sva_dfm_1,
      buf_acc_data_15_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_8_56_46_sva_dfm_1,
      buf_acc_data_15_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2478_nl = MUX_s_1_2_2(buf_acc_data_2_9_0_sva,
      buf_acc_data_2_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2478_nl,
      buf_acc_data_2_9_0_sva, or_dcpl_124);
  assign buf_acc_data_2_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_9_45_1_sva_dfm_1,
      buf_acc_data_2_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_9_56_46_sva_dfm_1,
      buf_acc_data_2_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2480_nl = MUX_s_1_2_2(buf_acc_data_15_7_0_sva,
      buf_acc_data_15_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2480_nl,
      buf_acc_data_15_7_0_sva, or_dcpl_124);
  assign buf_acc_data_15_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_7_45_1_sva_dfm_1,
      buf_acc_data_15_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_7_56_46_sva_dfm_1,
      buf_acc_data_15_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2482_nl = MUX_s_1_2_2(buf_acc_data_2_10_0_sva,
      buf_acc_data_2_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2482_nl,
      buf_acc_data_2_10_0_sva, or_dcpl_124);
  assign buf_acc_data_2_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_10_45_1_sva_dfm_1,
      buf_acc_data_2_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_10_56_46_sva_dfm_1,
      buf_acc_data_2_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2484_nl = MUX_s_1_2_2(buf_acc_data_15_6_0_sva,
      buf_acc_data_15_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2484_nl,
      buf_acc_data_15_6_0_sva, or_dcpl_124);
  assign buf_acc_data_15_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_6_45_1_sva_dfm_1,
      buf_acc_data_15_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_6_56_46_sva_dfm_1,
      buf_acc_data_15_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2486_nl = MUX_s_1_2_2(buf_acc_data_2_11_0_sva,
      buf_acc_data_2_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2486_nl,
      buf_acc_data_2_11_0_sva, or_dcpl_124);
  assign buf_acc_data_2_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_11_45_1_sva_dfm_1,
      buf_acc_data_2_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_11_56_46_sva_dfm_1,
      buf_acc_data_2_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2488_nl = MUX_s_1_2_2(buf_acc_data_15_5_0_sva,
      buf_acc_data_15_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2488_nl,
      buf_acc_data_15_5_0_sva, or_dcpl_124);
  assign buf_acc_data_15_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_5_45_1_sva_dfm_1,
      buf_acc_data_15_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_5_56_46_sva_dfm_1,
      buf_acc_data_15_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2490_nl = MUX_s_1_2_2(buf_acc_data_2_12_0_sva,
      buf_acc_data_2_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2490_nl,
      buf_acc_data_2_12_0_sva, or_dcpl_124);
  assign buf_acc_data_2_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_12_45_1_sva_dfm_1,
      buf_acc_data_2_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_12_56_46_sva_dfm_1,
      buf_acc_data_2_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2492_nl = MUX_s_1_2_2(buf_acc_data_15_4_0_sva,
      buf_acc_data_15_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2492_nl,
      buf_acc_data_15_4_0_sva, or_dcpl_124);
  assign buf_acc_data_15_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_4_45_1_sva_dfm_1,
      buf_acc_data_15_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_4_56_46_sva_dfm_1,
      buf_acc_data_15_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2494_nl = MUX_s_1_2_2(buf_acc_data_2_13_0_sva,
      buf_acc_data_2_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2494_nl,
      buf_acc_data_2_13_0_sva, or_dcpl_124);
  assign buf_acc_data_2_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_13_45_1_sva_dfm_1,
      buf_acc_data_2_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_13_56_46_sva_dfm_1,
      buf_acc_data_2_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2496_nl = MUX_s_1_2_2(buf_acc_data_15_3_0_sva,
      buf_acc_data_15_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2496_nl,
      buf_acc_data_15_3_0_sva, or_dcpl_124);
  assign buf_acc_data_15_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_3_45_1_sva_dfm_1,
      buf_acc_data_15_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_3_56_46_sva_dfm_1,
      buf_acc_data_15_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2498_nl = MUX_s_1_2_2(buf_acc_data_2_14_0_sva,
      buf_acc_data_2_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2498_nl,
      buf_acc_data_2_14_0_sva, or_dcpl_124);
  assign buf_acc_data_2_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_14_45_1_sva_dfm_1,
      buf_acc_data_2_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_14_56_46_sva_dfm_1,
      buf_acc_data_2_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2500_nl = MUX_s_1_2_2(buf_acc_data_15_2_0_sva,
      buf_acc_data_15_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2500_nl,
      buf_acc_data_15_2_0_sva, or_dcpl_124);
  assign buf_acc_data_15_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_2_45_1_sva_dfm_1,
      buf_acc_data_15_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_2_56_46_sva_dfm_1,
      buf_acc_data_15_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2502_nl = MUX_s_1_2_2(buf_acc_data_2_15_0_sva,
      buf_acc_data_2_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2502_nl,
      buf_acc_data_2_15_0_sva, or_dcpl_124);
  assign buf_acc_data_2_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_15_45_1_sva_dfm_1,
      buf_acc_data_2_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_15_56_46_sva_dfm_1,
      buf_acc_data_2_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2504_nl = MUX_s_1_2_2(buf_acc_data_15_1_0_sva,
      buf_acc_data_15_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2504_nl,
      buf_acc_data_15_1_0_sva, or_dcpl_124);
  assign buf_acc_data_15_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_1_45_1_sva_dfm_1,
      buf_acc_data_15_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_1_56_46_sva_dfm_1,
      buf_acc_data_15_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2506_nl = MUX_s_1_2_2(buf_acc_data_2_16_0_sva,
      buf_acc_data_2_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2506_nl,
      buf_acc_data_2_16_0_sva, or_dcpl_124);
  assign buf_acc_data_2_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_16_45_1_sva_dfm_1,
      buf_acc_data_2_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_16_56_46_sva_dfm_1,
      buf_acc_data_2_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2508_nl = MUX_s_1_2_2(buf_acc_data_15_0_0_sva,
      buf_acc_data_15_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_15_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2508_nl,
      buf_acc_data_15_0_0_sva, or_dcpl_124);
  assign buf_acc_data_15_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_15_0_45_1_sva_dfm_1,
      buf_acc_data_15_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_15_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_15_0_56_46_sva_dfm_1,
      buf_acc_data_15_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2510_nl = MUX_s_1_2_2(buf_acc_data_2_17_0_sva,
      buf_acc_data_2_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_2_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2510_nl,
      buf_acc_data_2_17_0_sva, or_dcpl_124);
  assign buf_acc_data_2_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_2_17_45_1_sva_dfm_1,
      buf_acc_data_2_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_2_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_2_17_56_46_sva_dfm_1,
      buf_acc_data_2_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2512_nl = MUX_s_1_2_2(buf_acc_data_14_17_0_sva,
      buf_acc_data_14_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2512_nl,
      buf_acc_data_14_17_0_sva, or_dcpl_124);
  assign buf_acc_data_14_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_17_45_1_sva_dfm_1,
      buf_acc_data_14_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_17_56_46_sva_dfm_1,
      buf_acc_data_14_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2514_nl = MUX_s_1_2_2(buf_acc_data_3_0_0_sva,
      buf_acc_data_3_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2514_nl,
      buf_acc_data_3_0_0_sva, or_dcpl_124);
  assign buf_acc_data_3_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_0_45_1_sva_dfm_1,
      buf_acc_data_3_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_0_56_46_sva_dfm_1,
      buf_acc_data_3_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2516_nl = MUX_s_1_2_2(buf_acc_data_14_16_0_sva,
      buf_acc_data_14_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2516_nl,
      buf_acc_data_14_16_0_sva, or_dcpl_124);
  assign buf_acc_data_14_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_16_45_1_sva_dfm_1,
      buf_acc_data_14_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_16_56_46_sva_dfm_1,
      buf_acc_data_14_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2518_nl = MUX_s_1_2_2(buf_acc_data_3_1_0_sva,
      buf_acc_data_3_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2518_nl,
      buf_acc_data_3_1_0_sva, or_dcpl_124);
  assign buf_acc_data_3_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_1_45_1_sva_dfm_1,
      buf_acc_data_3_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_1_56_46_sva_dfm_1,
      buf_acc_data_3_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2520_nl = MUX_s_1_2_2(buf_acc_data_14_15_0_sva,
      buf_acc_data_14_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2520_nl,
      buf_acc_data_14_15_0_sva, or_dcpl_124);
  assign buf_acc_data_14_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_15_45_1_sva_dfm_1,
      buf_acc_data_14_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_15_56_46_sva_dfm_1,
      buf_acc_data_14_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2522_nl = MUX_s_1_2_2(buf_acc_data_3_2_0_sva,
      buf_acc_data_3_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2522_nl,
      buf_acc_data_3_2_0_sva, or_dcpl_124);
  assign buf_acc_data_3_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_2_45_1_sva_dfm_1,
      buf_acc_data_3_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_2_56_46_sva_dfm_1,
      buf_acc_data_3_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2524_nl = MUX_s_1_2_2(buf_acc_data_14_14_0_sva,
      buf_acc_data_14_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2524_nl,
      buf_acc_data_14_14_0_sva, or_dcpl_124);
  assign buf_acc_data_14_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_14_45_1_sva_dfm_1,
      buf_acc_data_14_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_14_56_46_sva_dfm_1,
      buf_acc_data_14_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2526_nl = MUX_s_1_2_2(buf_acc_data_3_3_0_sva,
      buf_acc_data_3_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2526_nl,
      buf_acc_data_3_3_0_sva, or_dcpl_124);
  assign buf_acc_data_3_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_3_45_1_sva_dfm_1,
      buf_acc_data_3_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_3_56_46_sva_dfm_1,
      buf_acc_data_3_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2528_nl = MUX_s_1_2_2(buf_acc_data_14_13_0_sva,
      buf_acc_data_14_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2528_nl,
      buf_acc_data_14_13_0_sva, or_dcpl_124);
  assign buf_acc_data_14_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_13_45_1_sva_dfm_1,
      buf_acc_data_14_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_13_56_46_sva_dfm_1,
      buf_acc_data_14_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2530_nl = MUX_s_1_2_2(buf_acc_data_3_4_0_sva,
      buf_acc_data_3_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2530_nl,
      buf_acc_data_3_4_0_sva, or_dcpl_124);
  assign buf_acc_data_3_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_4_45_1_sva_dfm_1,
      buf_acc_data_3_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_4_56_46_sva_dfm_1,
      buf_acc_data_3_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2532_nl = MUX_s_1_2_2(buf_acc_data_14_12_0_sva,
      buf_acc_data_14_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2532_nl,
      buf_acc_data_14_12_0_sva, or_dcpl_124);
  assign buf_acc_data_14_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_12_45_1_sva_dfm_1,
      buf_acc_data_14_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_12_56_46_sva_dfm_1,
      buf_acc_data_14_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2534_nl = MUX_s_1_2_2(buf_acc_data_3_5_0_sva,
      buf_acc_data_3_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2534_nl,
      buf_acc_data_3_5_0_sva, or_dcpl_124);
  assign buf_acc_data_3_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_5_45_1_sva_dfm_1,
      buf_acc_data_3_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_5_56_46_sva_dfm_1,
      buf_acc_data_3_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2536_nl = MUX_s_1_2_2(buf_acc_data_14_11_0_sva,
      buf_acc_data_14_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2536_nl,
      buf_acc_data_14_11_0_sva, or_dcpl_124);
  assign buf_acc_data_14_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_11_45_1_sva_dfm_1,
      buf_acc_data_14_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_11_56_46_sva_dfm_1,
      buf_acc_data_14_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2538_nl = MUX_s_1_2_2(buf_acc_data_3_6_0_sva,
      buf_acc_data_3_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2538_nl,
      buf_acc_data_3_6_0_sva, or_dcpl_124);
  assign buf_acc_data_3_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_6_45_1_sva_dfm_1,
      buf_acc_data_3_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_6_56_46_sva_dfm_1,
      buf_acc_data_3_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2540_nl = MUX_s_1_2_2(buf_acc_data_14_10_0_sva,
      buf_acc_data_14_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2540_nl,
      buf_acc_data_14_10_0_sva, or_dcpl_124);
  assign buf_acc_data_14_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_10_45_1_sva_dfm_1,
      buf_acc_data_14_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_10_56_46_sva_dfm_1,
      buf_acc_data_14_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2542_nl = MUX_s_1_2_2(buf_acc_data_3_7_0_sva,
      buf_acc_data_3_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2542_nl,
      buf_acc_data_3_7_0_sva, or_dcpl_124);
  assign buf_acc_data_3_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_7_45_1_sva_dfm_1,
      buf_acc_data_3_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_7_56_46_sva_dfm_1,
      buf_acc_data_3_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2544_nl = MUX_s_1_2_2(buf_acc_data_14_9_0_sva,
      buf_acc_data_14_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2544_nl,
      buf_acc_data_14_9_0_sva, or_dcpl_124);
  assign buf_acc_data_14_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_9_45_1_sva_dfm_1,
      buf_acc_data_14_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_9_56_46_sva_dfm_1,
      buf_acc_data_14_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2546_nl = MUX_s_1_2_2(buf_acc_data_3_8_0_sva,
      buf_acc_data_3_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2546_nl,
      buf_acc_data_3_8_0_sva, or_dcpl_124);
  assign buf_acc_data_3_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_8_45_1_sva_dfm_1,
      buf_acc_data_3_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_8_56_46_sva_dfm_1,
      buf_acc_data_3_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2548_nl = MUX_s_1_2_2(buf_acc_data_14_8_0_sva,
      buf_acc_data_14_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2548_nl,
      buf_acc_data_14_8_0_sva, or_dcpl_124);
  assign buf_acc_data_14_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_8_45_1_sva_dfm_1,
      buf_acc_data_14_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_8_56_46_sva_dfm_1,
      buf_acc_data_14_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2550_nl = MUX_s_1_2_2(buf_acc_data_3_9_0_sva,
      buf_acc_data_3_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2550_nl,
      buf_acc_data_3_9_0_sva, or_dcpl_124);
  assign buf_acc_data_3_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_9_45_1_sva_dfm_1,
      buf_acc_data_3_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_9_56_46_sva_dfm_1,
      buf_acc_data_3_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2552_nl = MUX_s_1_2_2(buf_acc_data_14_7_0_sva,
      buf_acc_data_14_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2552_nl,
      buf_acc_data_14_7_0_sva, or_dcpl_124);
  assign buf_acc_data_14_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_7_45_1_sva_dfm_1,
      buf_acc_data_14_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_7_56_46_sva_dfm_1,
      buf_acc_data_14_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2554_nl = MUX_s_1_2_2(buf_acc_data_3_10_0_sva,
      buf_acc_data_3_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2554_nl,
      buf_acc_data_3_10_0_sva, or_dcpl_124);
  assign buf_acc_data_3_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_10_45_1_sva_dfm_1,
      buf_acc_data_3_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_10_56_46_sva_dfm_1,
      buf_acc_data_3_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2556_nl = MUX_s_1_2_2(buf_acc_data_14_6_0_sva,
      buf_acc_data_14_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2556_nl,
      buf_acc_data_14_6_0_sva, or_dcpl_124);
  assign buf_acc_data_14_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_6_45_1_sva_dfm_1,
      buf_acc_data_14_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_6_56_46_sva_dfm_1,
      buf_acc_data_14_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2558_nl = MUX_s_1_2_2(buf_acc_data_3_11_0_sva,
      buf_acc_data_3_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2558_nl,
      buf_acc_data_3_11_0_sva, or_dcpl_124);
  assign buf_acc_data_3_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_11_45_1_sva_dfm_1,
      buf_acc_data_3_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_11_56_46_sva_dfm_1,
      buf_acc_data_3_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2560_nl = MUX_s_1_2_2(buf_acc_data_14_5_0_sva,
      buf_acc_data_14_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2560_nl,
      buf_acc_data_14_5_0_sva, or_dcpl_124);
  assign buf_acc_data_14_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_5_45_1_sva_dfm_1,
      buf_acc_data_14_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_5_56_46_sva_dfm_1,
      buf_acc_data_14_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2562_nl = MUX_s_1_2_2(buf_acc_data_3_12_0_sva,
      buf_acc_data_3_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2562_nl,
      buf_acc_data_3_12_0_sva, or_dcpl_124);
  assign buf_acc_data_3_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_12_45_1_sva_dfm_1,
      buf_acc_data_3_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_12_56_46_sva_dfm_1,
      buf_acc_data_3_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2564_nl = MUX_s_1_2_2(buf_acc_data_14_4_0_sva,
      buf_acc_data_14_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2564_nl,
      buf_acc_data_14_4_0_sva, or_dcpl_124);
  assign buf_acc_data_14_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_4_45_1_sva_dfm_1,
      buf_acc_data_14_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_4_56_46_sva_dfm_1,
      buf_acc_data_14_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2566_nl = MUX_s_1_2_2(buf_acc_data_3_13_0_sva,
      buf_acc_data_3_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2566_nl,
      buf_acc_data_3_13_0_sva, or_dcpl_124);
  assign buf_acc_data_3_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_13_45_1_sva_dfm_1,
      buf_acc_data_3_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_13_56_46_sva_dfm_1,
      buf_acc_data_3_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2568_nl = MUX_s_1_2_2(buf_acc_data_14_3_0_sva,
      buf_acc_data_14_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2568_nl,
      buf_acc_data_14_3_0_sva, or_dcpl_124);
  assign buf_acc_data_14_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_3_45_1_sva_dfm_1,
      buf_acc_data_14_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_3_56_46_sva_dfm_1,
      buf_acc_data_14_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2570_nl = MUX_s_1_2_2(buf_acc_data_3_14_0_sva,
      buf_acc_data_3_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2570_nl,
      buf_acc_data_3_14_0_sva, or_dcpl_124);
  assign buf_acc_data_3_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_14_45_1_sva_dfm_1,
      buf_acc_data_3_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_14_56_46_sva_dfm_1,
      buf_acc_data_3_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2572_nl = MUX_s_1_2_2(buf_acc_data_14_2_0_sva,
      buf_acc_data_14_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2572_nl,
      buf_acc_data_14_2_0_sva, or_dcpl_124);
  assign buf_acc_data_14_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_2_45_1_sva_dfm_1,
      buf_acc_data_14_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_2_56_46_sva_dfm_1,
      buf_acc_data_14_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2574_nl = MUX_s_1_2_2(buf_acc_data_3_15_0_sva,
      buf_acc_data_3_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2574_nl,
      buf_acc_data_3_15_0_sva, or_dcpl_124);
  assign buf_acc_data_3_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_15_45_1_sva_dfm_1,
      buf_acc_data_3_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_15_56_46_sva_dfm_1,
      buf_acc_data_3_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2576_nl = MUX_s_1_2_2(buf_acc_data_14_1_0_sva,
      buf_acc_data_14_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2576_nl,
      buf_acc_data_14_1_0_sva, or_dcpl_124);
  assign buf_acc_data_14_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_1_45_1_sva_dfm_1,
      buf_acc_data_14_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_1_56_46_sva_dfm_1,
      buf_acc_data_14_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2578_nl = MUX_s_1_2_2(buf_acc_data_3_16_0_sva,
      buf_acc_data_3_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2578_nl,
      buf_acc_data_3_16_0_sva, or_dcpl_124);
  assign buf_acc_data_3_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_16_45_1_sva_dfm_1,
      buf_acc_data_3_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_16_56_46_sva_dfm_1,
      buf_acc_data_3_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2580_nl = MUX_s_1_2_2(buf_acc_data_14_0_0_sva,
      buf_acc_data_14_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_14_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2580_nl,
      buf_acc_data_14_0_0_sva, or_dcpl_124);
  assign buf_acc_data_14_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_14_0_45_1_sva_dfm_1,
      buf_acc_data_14_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_14_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_14_0_56_46_sva_dfm_1,
      buf_acc_data_14_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2582_nl = MUX_s_1_2_2(buf_acc_data_3_17_0_sva,
      buf_acc_data_3_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_3_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2582_nl,
      buf_acc_data_3_17_0_sva, or_dcpl_124);
  assign buf_acc_data_3_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_3_17_45_1_sva_dfm_1,
      buf_acc_data_3_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_3_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_3_17_56_46_sva_dfm_1,
      buf_acc_data_3_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2584_nl = MUX_s_1_2_2(buf_acc_data_13_17_0_sva,
      buf_acc_data_13_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2584_nl,
      buf_acc_data_13_17_0_sva, or_dcpl_124);
  assign buf_acc_data_13_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_17_45_1_sva_dfm_1,
      buf_acc_data_13_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_17_56_46_sva_dfm_1,
      buf_acc_data_13_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2586_nl = MUX_s_1_2_2(buf_acc_data_4_0_0_sva,
      buf_acc_data_4_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2586_nl,
      buf_acc_data_4_0_0_sva, or_dcpl_124);
  assign buf_acc_data_4_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_0_45_1_sva_dfm_1,
      buf_acc_data_4_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_0_56_46_sva_dfm_1,
      buf_acc_data_4_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2588_nl = MUX_s_1_2_2(buf_acc_data_13_16_0_sva,
      buf_acc_data_13_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2588_nl,
      buf_acc_data_13_16_0_sva, or_dcpl_124);
  assign buf_acc_data_13_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_16_45_1_sva_dfm_1,
      buf_acc_data_13_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_16_56_46_sva_dfm_1,
      buf_acc_data_13_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2590_nl = MUX_s_1_2_2(buf_acc_data_4_1_0_sva,
      buf_acc_data_4_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2590_nl,
      buf_acc_data_4_1_0_sva, or_dcpl_124);
  assign buf_acc_data_4_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_1_45_1_sva_dfm_1,
      buf_acc_data_4_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_1_56_46_sva_dfm_1,
      buf_acc_data_4_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2592_nl = MUX_s_1_2_2(buf_acc_data_13_15_0_sva,
      buf_acc_data_13_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2592_nl,
      buf_acc_data_13_15_0_sva, or_dcpl_124);
  assign buf_acc_data_13_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_15_45_1_sva_dfm_1,
      buf_acc_data_13_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_15_56_46_sva_dfm_1,
      buf_acc_data_13_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2594_nl = MUX_s_1_2_2(buf_acc_data_4_2_0_sva,
      buf_acc_data_4_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2594_nl,
      buf_acc_data_4_2_0_sva, or_dcpl_124);
  assign buf_acc_data_4_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_2_45_1_sva_dfm_1,
      buf_acc_data_4_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_2_56_46_sva_dfm_1,
      buf_acc_data_4_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2596_nl = MUX_s_1_2_2(buf_acc_data_13_14_0_sva,
      buf_acc_data_13_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2596_nl,
      buf_acc_data_13_14_0_sva, or_dcpl_124);
  assign buf_acc_data_13_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_14_45_1_sva_dfm_1,
      buf_acc_data_13_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_14_56_46_sva_dfm_1,
      buf_acc_data_13_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2598_nl = MUX_s_1_2_2(buf_acc_data_4_3_0_sva,
      buf_acc_data_4_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2598_nl,
      buf_acc_data_4_3_0_sva, or_dcpl_124);
  assign buf_acc_data_4_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_3_45_1_sva_dfm_1,
      buf_acc_data_4_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_3_56_46_sva_dfm_1,
      buf_acc_data_4_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2600_nl = MUX_s_1_2_2(buf_acc_data_13_13_0_sva,
      buf_acc_data_13_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2600_nl,
      buf_acc_data_13_13_0_sva, or_dcpl_124);
  assign buf_acc_data_13_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_13_45_1_sva_dfm_1,
      buf_acc_data_13_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_13_56_46_sva_dfm_1,
      buf_acc_data_13_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2602_nl = MUX_s_1_2_2(buf_acc_data_4_4_0_sva,
      buf_acc_data_4_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2602_nl,
      buf_acc_data_4_4_0_sva, or_dcpl_124);
  assign buf_acc_data_4_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_4_45_1_sva_dfm_1,
      buf_acc_data_4_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_4_56_46_sva_dfm_1,
      buf_acc_data_4_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2604_nl = MUX_s_1_2_2(buf_acc_data_13_12_0_sva,
      buf_acc_data_13_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2604_nl,
      buf_acc_data_13_12_0_sva, or_dcpl_124);
  assign buf_acc_data_13_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_12_45_1_sva_dfm_1,
      buf_acc_data_13_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_12_56_46_sva_dfm_1,
      buf_acc_data_13_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2606_nl = MUX_s_1_2_2(buf_acc_data_4_5_0_sva,
      buf_acc_data_4_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2606_nl,
      buf_acc_data_4_5_0_sva, or_dcpl_124);
  assign buf_acc_data_4_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_5_45_1_sva_dfm_1,
      buf_acc_data_4_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_5_56_46_sva_dfm_1,
      buf_acc_data_4_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2608_nl = MUX_s_1_2_2(buf_acc_data_13_11_0_sva,
      buf_acc_data_13_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2608_nl,
      buf_acc_data_13_11_0_sva, or_dcpl_124);
  assign buf_acc_data_13_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_11_45_1_sva_dfm_1,
      buf_acc_data_13_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_11_56_46_sva_dfm_1,
      buf_acc_data_13_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2610_nl = MUX_s_1_2_2(buf_acc_data_4_6_0_sva,
      buf_acc_data_4_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2610_nl,
      buf_acc_data_4_6_0_sva, or_dcpl_124);
  assign buf_acc_data_4_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_6_45_1_sva_dfm_1,
      buf_acc_data_4_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_6_56_46_sva_dfm_1,
      buf_acc_data_4_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2612_nl = MUX_s_1_2_2(buf_acc_data_13_10_0_sva,
      buf_acc_data_13_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2612_nl,
      buf_acc_data_13_10_0_sva, or_dcpl_124);
  assign buf_acc_data_13_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_10_45_1_sva_dfm_1,
      buf_acc_data_13_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_10_56_46_sva_dfm_1,
      buf_acc_data_13_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2614_nl = MUX_s_1_2_2(buf_acc_data_4_7_0_sva,
      buf_acc_data_4_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2614_nl,
      buf_acc_data_4_7_0_sva, or_dcpl_124);
  assign buf_acc_data_4_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_7_45_1_sva_dfm_1,
      buf_acc_data_4_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_7_56_46_sva_dfm_1,
      buf_acc_data_4_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2616_nl = MUX_s_1_2_2(buf_acc_data_13_9_0_sva,
      buf_acc_data_13_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2616_nl,
      buf_acc_data_13_9_0_sva, or_dcpl_124);
  assign buf_acc_data_13_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_9_45_1_sva_dfm_1,
      buf_acc_data_13_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_9_56_46_sva_dfm_1,
      buf_acc_data_13_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2618_nl = MUX_s_1_2_2(buf_acc_data_4_8_0_sva,
      buf_acc_data_4_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2618_nl,
      buf_acc_data_4_8_0_sva, or_dcpl_124);
  assign buf_acc_data_4_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_8_45_1_sva_dfm_1,
      buf_acc_data_4_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_8_56_46_sva_dfm_1,
      buf_acc_data_4_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2620_nl = MUX_s_1_2_2(buf_acc_data_13_8_0_sva,
      buf_acc_data_13_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2620_nl,
      buf_acc_data_13_8_0_sva, or_dcpl_124);
  assign buf_acc_data_13_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_8_45_1_sva_dfm_1,
      buf_acc_data_13_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_8_56_46_sva_dfm_1,
      buf_acc_data_13_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2622_nl = MUX_s_1_2_2(buf_acc_data_4_9_0_sva,
      buf_acc_data_4_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2622_nl,
      buf_acc_data_4_9_0_sva, or_dcpl_124);
  assign buf_acc_data_4_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_9_45_1_sva_dfm_1,
      buf_acc_data_4_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_9_56_46_sva_dfm_1,
      buf_acc_data_4_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2624_nl = MUX_s_1_2_2(buf_acc_data_13_7_0_sva,
      buf_acc_data_13_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2624_nl,
      buf_acc_data_13_7_0_sva, or_dcpl_124);
  assign buf_acc_data_13_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_7_45_1_sva_dfm_1,
      buf_acc_data_13_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_7_56_46_sva_dfm_1,
      buf_acc_data_13_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2626_nl = MUX_s_1_2_2(buf_acc_data_4_10_0_sva,
      buf_acc_data_4_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2626_nl,
      buf_acc_data_4_10_0_sva, or_dcpl_124);
  assign buf_acc_data_4_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_10_45_1_sva_dfm_1,
      buf_acc_data_4_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_10_56_46_sva_dfm_1,
      buf_acc_data_4_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2628_nl = MUX_s_1_2_2(buf_acc_data_13_6_0_sva,
      buf_acc_data_13_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2628_nl,
      buf_acc_data_13_6_0_sva, or_dcpl_124);
  assign buf_acc_data_13_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_6_45_1_sva_dfm_1,
      buf_acc_data_13_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_6_56_46_sva_dfm_1,
      buf_acc_data_13_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2630_nl = MUX_s_1_2_2(buf_acc_data_4_11_0_sva,
      buf_acc_data_4_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2630_nl,
      buf_acc_data_4_11_0_sva, or_dcpl_124);
  assign buf_acc_data_4_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_11_45_1_sva_dfm_1,
      buf_acc_data_4_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_11_56_46_sva_dfm_1,
      buf_acc_data_4_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2632_nl = MUX_s_1_2_2(buf_acc_data_13_5_0_sva,
      buf_acc_data_13_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2632_nl,
      buf_acc_data_13_5_0_sva, or_dcpl_124);
  assign buf_acc_data_13_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_5_45_1_sva_dfm_1,
      buf_acc_data_13_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_5_56_46_sva_dfm_1,
      buf_acc_data_13_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2634_nl = MUX_s_1_2_2(buf_acc_data_4_12_0_sva,
      buf_acc_data_4_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2634_nl,
      buf_acc_data_4_12_0_sva, or_dcpl_124);
  assign buf_acc_data_4_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_12_45_1_sva_dfm_1,
      buf_acc_data_4_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_12_56_46_sva_dfm_1,
      buf_acc_data_4_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2636_nl = MUX_s_1_2_2(buf_acc_data_13_4_0_sva,
      buf_acc_data_13_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2636_nl,
      buf_acc_data_13_4_0_sva, or_dcpl_124);
  assign buf_acc_data_13_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_4_45_1_sva_dfm_1,
      buf_acc_data_13_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_4_56_46_sva_dfm_1,
      buf_acc_data_13_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2638_nl = MUX_s_1_2_2(buf_acc_data_4_13_0_sva,
      buf_acc_data_4_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2638_nl,
      buf_acc_data_4_13_0_sva, or_dcpl_124);
  assign buf_acc_data_4_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_13_45_1_sva_dfm_1,
      buf_acc_data_4_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_13_56_46_sva_dfm_1,
      buf_acc_data_4_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2640_nl = MUX_s_1_2_2(buf_acc_data_13_3_0_sva,
      buf_acc_data_13_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2640_nl,
      buf_acc_data_13_3_0_sva, or_dcpl_124);
  assign buf_acc_data_13_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_3_45_1_sva_dfm_1,
      buf_acc_data_13_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_3_56_46_sva_dfm_1,
      buf_acc_data_13_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2642_nl = MUX_s_1_2_2(buf_acc_data_4_14_0_sva,
      buf_acc_data_4_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2642_nl,
      buf_acc_data_4_14_0_sva, or_dcpl_124);
  assign buf_acc_data_4_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_14_45_1_sva_dfm_1,
      buf_acc_data_4_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_14_56_46_sva_dfm_1,
      buf_acc_data_4_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2644_nl = MUX_s_1_2_2(buf_acc_data_13_2_0_sva,
      buf_acc_data_13_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2644_nl,
      buf_acc_data_13_2_0_sva, or_dcpl_124);
  assign buf_acc_data_13_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_2_45_1_sva_dfm_1,
      buf_acc_data_13_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_2_56_46_sva_dfm_1,
      buf_acc_data_13_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2646_nl = MUX_s_1_2_2(buf_acc_data_4_15_0_sva,
      buf_acc_data_4_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2646_nl,
      buf_acc_data_4_15_0_sva, or_dcpl_124);
  assign buf_acc_data_4_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_15_45_1_sva_dfm_1,
      buf_acc_data_4_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_15_56_46_sva_dfm_1,
      buf_acc_data_4_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2648_nl = MUX_s_1_2_2(buf_acc_data_13_1_0_sva,
      buf_acc_data_13_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2648_nl,
      buf_acc_data_13_1_0_sva, or_dcpl_124);
  assign buf_acc_data_13_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_1_45_1_sva_dfm_1,
      buf_acc_data_13_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_1_56_46_sva_dfm_1,
      buf_acc_data_13_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2650_nl = MUX_s_1_2_2(buf_acc_data_4_16_0_sva,
      buf_acc_data_4_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2650_nl,
      buf_acc_data_4_16_0_sva, or_dcpl_124);
  assign buf_acc_data_4_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_16_45_1_sva_dfm_1,
      buf_acc_data_4_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_16_56_46_sva_dfm_1,
      buf_acc_data_4_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2652_nl = MUX_s_1_2_2(buf_acc_data_13_0_0_sva,
      buf_acc_data_13_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_13_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2652_nl,
      buf_acc_data_13_0_0_sva, or_dcpl_124);
  assign buf_acc_data_13_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_13_0_45_1_sva_dfm_1,
      buf_acc_data_13_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_13_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_13_0_56_46_sva_dfm_1,
      buf_acc_data_13_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2654_nl = MUX_s_1_2_2(buf_acc_data_4_17_0_sva,
      buf_acc_data_4_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_4_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2654_nl,
      buf_acc_data_4_17_0_sva, or_dcpl_124);
  assign buf_acc_data_4_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_4_17_45_1_sva_dfm_1,
      buf_acc_data_4_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_4_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_4_17_56_46_sva_dfm_1,
      buf_acc_data_4_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2656_nl = MUX_s_1_2_2(buf_acc_data_12_17_0_sva,
      buf_acc_data_12_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2656_nl,
      buf_acc_data_12_17_0_sva, or_dcpl_124);
  assign buf_acc_data_12_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_17_45_1_sva_dfm_1,
      buf_acc_data_12_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_17_56_46_sva_dfm_1,
      buf_acc_data_12_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2658_nl = MUX_s_1_2_2(buf_acc_data_5_0_0_sva,
      buf_acc_data_5_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2658_nl,
      buf_acc_data_5_0_0_sva, or_dcpl_124);
  assign buf_acc_data_5_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_0_45_1_sva_dfm_1,
      buf_acc_data_5_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_0_56_46_sva_dfm_1,
      buf_acc_data_5_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2660_nl = MUX_s_1_2_2(buf_acc_data_12_16_0_sva,
      buf_acc_data_12_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2660_nl,
      buf_acc_data_12_16_0_sva, or_dcpl_124);
  assign buf_acc_data_12_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_16_45_1_sva_dfm_1,
      buf_acc_data_12_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_16_56_46_sva_dfm_1,
      buf_acc_data_12_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2662_nl = MUX_s_1_2_2(buf_acc_data_5_1_0_sva,
      buf_acc_data_5_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2662_nl,
      buf_acc_data_5_1_0_sva, or_dcpl_124);
  assign buf_acc_data_5_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_1_45_1_sva_dfm_1,
      buf_acc_data_5_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_1_56_46_sva_dfm_1,
      buf_acc_data_5_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2664_nl = MUX_s_1_2_2(buf_acc_data_12_15_0_sva,
      buf_acc_data_12_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2664_nl,
      buf_acc_data_12_15_0_sva, or_dcpl_124);
  assign buf_acc_data_12_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_15_45_1_sva_dfm_1,
      buf_acc_data_12_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_15_56_46_sva_dfm_1,
      buf_acc_data_12_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2666_nl = MUX_s_1_2_2(buf_acc_data_5_2_0_sva,
      buf_acc_data_5_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2666_nl,
      buf_acc_data_5_2_0_sva, or_dcpl_124);
  assign buf_acc_data_5_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_2_45_1_sva_dfm_1,
      buf_acc_data_5_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_2_56_46_sva_dfm_1,
      buf_acc_data_5_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2668_nl = MUX_s_1_2_2(buf_acc_data_12_14_0_sva,
      buf_acc_data_12_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2668_nl,
      buf_acc_data_12_14_0_sva, or_dcpl_124);
  assign buf_acc_data_12_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_14_45_1_sva_dfm_1,
      buf_acc_data_12_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_14_56_46_sva_dfm_1,
      buf_acc_data_12_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2670_nl = MUX_s_1_2_2(buf_acc_data_5_3_0_sva,
      buf_acc_data_5_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2670_nl,
      buf_acc_data_5_3_0_sva, or_dcpl_124);
  assign buf_acc_data_5_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_3_45_1_sva_dfm_1,
      buf_acc_data_5_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_3_56_46_sva_dfm_1,
      buf_acc_data_5_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2672_nl = MUX_s_1_2_2(buf_acc_data_12_13_0_sva,
      buf_acc_data_12_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2672_nl,
      buf_acc_data_12_13_0_sva, or_dcpl_124);
  assign buf_acc_data_12_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_13_45_1_sva_dfm_1,
      buf_acc_data_12_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_13_56_46_sva_dfm_1,
      buf_acc_data_12_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2674_nl = MUX_s_1_2_2(buf_acc_data_5_4_0_sva,
      buf_acc_data_5_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2674_nl,
      buf_acc_data_5_4_0_sva, or_dcpl_124);
  assign buf_acc_data_5_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_4_45_1_sva_dfm_1,
      buf_acc_data_5_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_4_56_46_sva_dfm_1,
      buf_acc_data_5_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2676_nl = MUX_s_1_2_2(buf_acc_data_12_12_0_sva,
      buf_acc_data_12_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2676_nl,
      buf_acc_data_12_12_0_sva, or_dcpl_124);
  assign buf_acc_data_12_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_12_45_1_sva_dfm_1,
      buf_acc_data_12_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_12_56_46_sva_dfm_1,
      buf_acc_data_12_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2678_nl = MUX_s_1_2_2(buf_acc_data_5_5_0_sva,
      buf_acc_data_5_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2678_nl,
      buf_acc_data_5_5_0_sva, or_dcpl_124);
  assign buf_acc_data_5_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_5_45_1_sva_dfm_1,
      buf_acc_data_5_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_5_56_46_sva_dfm_1,
      buf_acc_data_5_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2680_nl = MUX_s_1_2_2(buf_acc_data_12_11_0_sva,
      buf_acc_data_12_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2680_nl,
      buf_acc_data_12_11_0_sva, or_dcpl_124);
  assign buf_acc_data_12_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_11_45_1_sva_dfm_1,
      buf_acc_data_12_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_11_56_46_sva_dfm_1,
      buf_acc_data_12_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2682_nl = MUX_s_1_2_2(buf_acc_data_5_6_0_sva,
      buf_acc_data_5_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2682_nl,
      buf_acc_data_5_6_0_sva, or_dcpl_124);
  assign buf_acc_data_5_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_6_45_1_sva_dfm_1,
      buf_acc_data_5_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_6_56_46_sva_dfm_1,
      buf_acc_data_5_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2684_nl = MUX_s_1_2_2(buf_acc_data_12_10_0_sva,
      buf_acc_data_12_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2684_nl,
      buf_acc_data_12_10_0_sva, or_dcpl_124);
  assign buf_acc_data_12_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_10_45_1_sva_dfm_1,
      buf_acc_data_12_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_10_56_46_sva_dfm_1,
      buf_acc_data_12_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2686_nl = MUX_s_1_2_2(buf_acc_data_5_7_0_sva,
      buf_acc_data_5_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2686_nl,
      buf_acc_data_5_7_0_sva, or_dcpl_124);
  assign buf_acc_data_5_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_7_45_1_sva_dfm_1,
      buf_acc_data_5_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_7_56_46_sva_dfm_1,
      buf_acc_data_5_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2688_nl = MUX_s_1_2_2(buf_acc_data_12_9_0_sva,
      buf_acc_data_12_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2688_nl,
      buf_acc_data_12_9_0_sva, or_dcpl_124);
  assign buf_acc_data_12_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_9_45_1_sva_dfm_1,
      buf_acc_data_12_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_9_56_46_sva_dfm_1,
      buf_acc_data_12_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2690_nl = MUX_s_1_2_2(buf_acc_data_5_8_0_sva,
      buf_acc_data_5_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2690_nl,
      buf_acc_data_5_8_0_sva, or_dcpl_124);
  assign buf_acc_data_5_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_8_45_1_sva_dfm_1,
      buf_acc_data_5_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_8_56_46_sva_dfm_1,
      buf_acc_data_5_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2692_nl = MUX_s_1_2_2(buf_acc_data_12_8_0_sva,
      buf_acc_data_12_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2692_nl,
      buf_acc_data_12_8_0_sva, or_dcpl_124);
  assign buf_acc_data_12_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_8_45_1_sva_dfm_1,
      buf_acc_data_12_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_8_56_46_sva_dfm_1,
      buf_acc_data_12_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2694_nl = MUX_s_1_2_2(buf_acc_data_5_9_0_sva,
      buf_acc_data_5_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2694_nl,
      buf_acc_data_5_9_0_sva, or_dcpl_124);
  assign buf_acc_data_5_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_9_45_1_sva_dfm_1,
      buf_acc_data_5_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_9_56_46_sva_dfm_1,
      buf_acc_data_5_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2696_nl = MUX_s_1_2_2(buf_acc_data_12_7_0_sva,
      buf_acc_data_12_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2696_nl,
      buf_acc_data_12_7_0_sva, or_dcpl_124);
  assign buf_acc_data_12_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_7_45_1_sva_dfm_1,
      buf_acc_data_12_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_7_56_46_sva_dfm_1,
      buf_acc_data_12_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2698_nl = MUX_s_1_2_2(buf_acc_data_5_10_0_sva,
      buf_acc_data_5_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2698_nl,
      buf_acc_data_5_10_0_sva, or_dcpl_124);
  assign buf_acc_data_5_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_10_45_1_sva_dfm_1,
      buf_acc_data_5_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_10_56_46_sva_dfm_1,
      buf_acc_data_5_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2700_nl = MUX_s_1_2_2(buf_acc_data_12_6_0_sva,
      buf_acc_data_12_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2700_nl,
      buf_acc_data_12_6_0_sva, or_dcpl_124);
  assign buf_acc_data_12_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_6_45_1_sva_dfm_1,
      buf_acc_data_12_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_6_56_46_sva_dfm_1,
      buf_acc_data_12_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2702_nl = MUX_s_1_2_2(buf_acc_data_5_11_0_sva,
      buf_acc_data_5_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2702_nl,
      buf_acc_data_5_11_0_sva, or_dcpl_124);
  assign buf_acc_data_5_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_11_45_1_sva_dfm_1,
      buf_acc_data_5_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_11_56_46_sva_dfm_1,
      buf_acc_data_5_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2704_nl = MUX_s_1_2_2(buf_acc_data_12_5_0_sva,
      buf_acc_data_12_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2704_nl,
      buf_acc_data_12_5_0_sva, or_dcpl_124);
  assign buf_acc_data_12_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_5_45_1_sva_dfm_1,
      buf_acc_data_12_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_5_56_46_sva_dfm_1,
      buf_acc_data_12_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2706_nl = MUX_s_1_2_2(buf_acc_data_5_12_0_sva,
      buf_acc_data_5_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2706_nl,
      buf_acc_data_5_12_0_sva, or_dcpl_124);
  assign buf_acc_data_5_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_12_45_1_sva_dfm_1,
      buf_acc_data_5_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_12_56_46_sva_dfm_1,
      buf_acc_data_5_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2708_nl = MUX_s_1_2_2(buf_acc_data_12_4_0_sva,
      buf_acc_data_12_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2708_nl,
      buf_acc_data_12_4_0_sva, or_dcpl_124);
  assign buf_acc_data_12_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_4_45_1_sva_dfm_1,
      buf_acc_data_12_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_4_56_46_sva_dfm_1,
      buf_acc_data_12_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2710_nl = MUX_s_1_2_2(buf_acc_data_5_13_0_sva,
      buf_acc_data_5_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2710_nl,
      buf_acc_data_5_13_0_sva, or_dcpl_124);
  assign buf_acc_data_5_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_13_45_1_sva_dfm_1,
      buf_acc_data_5_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_13_56_46_sva_dfm_1,
      buf_acc_data_5_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2712_nl = MUX_s_1_2_2(buf_acc_data_12_3_0_sva,
      buf_acc_data_12_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2712_nl,
      buf_acc_data_12_3_0_sva, or_dcpl_124);
  assign buf_acc_data_12_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_3_45_1_sva_dfm_1,
      buf_acc_data_12_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_3_56_46_sva_dfm_1,
      buf_acc_data_12_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2714_nl = MUX_s_1_2_2(buf_acc_data_5_14_0_sva,
      buf_acc_data_5_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2714_nl,
      buf_acc_data_5_14_0_sva, or_dcpl_124);
  assign buf_acc_data_5_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_14_45_1_sva_dfm_1,
      buf_acc_data_5_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_14_56_46_sva_dfm_1,
      buf_acc_data_5_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2716_nl = MUX_s_1_2_2(buf_acc_data_12_2_0_sva,
      buf_acc_data_12_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2716_nl,
      buf_acc_data_12_2_0_sva, or_dcpl_124);
  assign buf_acc_data_12_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_2_45_1_sva_dfm_1,
      buf_acc_data_12_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_2_56_46_sva_dfm_1,
      buf_acc_data_12_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2718_nl = MUX_s_1_2_2(buf_acc_data_5_15_0_sva,
      buf_acc_data_5_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2718_nl,
      buf_acc_data_5_15_0_sva, or_dcpl_124);
  assign buf_acc_data_5_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_15_45_1_sva_dfm_1,
      buf_acc_data_5_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_15_56_46_sva_dfm_1,
      buf_acc_data_5_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2720_nl = MUX_s_1_2_2(buf_acc_data_12_1_0_sva,
      buf_acc_data_12_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2720_nl,
      buf_acc_data_12_1_0_sva, or_dcpl_124);
  assign buf_acc_data_12_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_1_45_1_sva_dfm_1,
      buf_acc_data_12_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_1_56_46_sva_dfm_1,
      buf_acc_data_12_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2722_nl = MUX_s_1_2_2(buf_acc_data_5_16_0_sva,
      buf_acc_data_5_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2722_nl,
      buf_acc_data_5_16_0_sva, or_dcpl_124);
  assign buf_acc_data_5_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_16_45_1_sva_dfm_1,
      buf_acc_data_5_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_16_56_46_sva_dfm_1,
      buf_acc_data_5_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2724_nl = MUX_s_1_2_2(buf_acc_data_12_0_0_sva,
      buf_acc_data_12_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_12_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2724_nl,
      buf_acc_data_12_0_0_sva, or_dcpl_124);
  assign buf_acc_data_12_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_12_0_45_1_sva_dfm_1,
      buf_acc_data_12_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_12_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_12_0_56_46_sva_dfm_1,
      buf_acc_data_12_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2726_nl = MUX_s_1_2_2(buf_acc_data_5_17_0_sva,
      buf_acc_data_5_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_5_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2726_nl,
      buf_acc_data_5_17_0_sva, or_dcpl_124);
  assign buf_acc_data_5_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_5_17_45_1_sva_dfm_1,
      buf_acc_data_5_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_5_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_5_17_56_46_sva_dfm_1,
      buf_acc_data_5_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2728_nl = MUX_s_1_2_2(buf_acc_data_11_17_0_sva,
      buf_acc_data_11_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2728_nl,
      buf_acc_data_11_17_0_sva, or_dcpl_124);
  assign buf_acc_data_11_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_17_45_1_sva_dfm_1,
      buf_acc_data_11_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_17_56_46_sva_dfm_1,
      buf_acc_data_11_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2730_nl = MUX_s_1_2_2(buf_acc_data_6_0_0_sva,
      buf_acc_data_6_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2730_nl,
      buf_acc_data_6_0_0_sva, or_dcpl_124);
  assign buf_acc_data_6_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_0_45_1_sva_dfm_1,
      buf_acc_data_6_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_0_56_46_sva_dfm_1,
      buf_acc_data_6_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2732_nl = MUX_s_1_2_2(buf_acc_data_11_16_0_sva,
      buf_acc_data_11_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2732_nl,
      buf_acc_data_11_16_0_sva, or_dcpl_124);
  assign buf_acc_data_11_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_16_45_1_sva_dfm_1,
      buf_acc_data_11_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_16_56_46_sva_dfm_1,
      buf_acc_data_11_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2734_nl = MUX_s_1_2_2(buf_acc_data_6_1_0_sva,
      buf_acc_data_6_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2734_nl,
      buf_acc_data_6_1_0_sva, or_dcpl_124);
  assign buf_acc_data_6_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_1_45_1_sva_dfm_1,
      buf_acc_data_6_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_1_56_46_sva_dfm_1,
      buf_acc_data_6_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2736_nl = MUX_s_1_2_2(buf_acc_data_11_15_0_sva,
      buf_acc_data_11_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2736_nl,
      buf_acc_data_11_15_0_sva, or_dcpl_124);
  assign buf_acc_data_11_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_15_45_1_sva_dfm_1,
      buf_acc_data_11_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_15_56_46_sva_dfm_1,
      buf_acc_data_11_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2738_nl = MUX_s_1_2_2(buf_acc_data_6_2_0_sva,
      buf_acc_data_6_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2738_nl,
      buf_acc_data_6_2_0_sva, or_dcpl_124);
  assign buf_acc_data_6_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_2_45_1_sva_dfm_1,
      buf_acc_data_6_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_2_56_46_sva_dfm_1,
      buf_acc_data_6_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2740_nl = MUX_s_1_2_2(buf_acc_data_11_14_0_sva,
      buf_acc_data_11_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2740_nl,
      buf_acc_data_11_14_0_sva, or_dcpl_124);
  assign buf_acc_data_11_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_14_45_1_sva_dfm_1,
      buf_acc_data_11_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_14_56_46_sva_dfm_1,
      buf_acc_data_11_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2742_nl = MUX_s_1_2_2(buf_acc_data_6_3_0_sva,
      buf_acc_data_6_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2742_nl,
      buf_acc_data_6_3_0_sva, or_dcpl_124);
  assign buf_acc_data_6_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_3_45_1_sva_dfm_1,
      buf_acc_data_6_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_3_56_46_sva_dfm_1,
      buf_acc_data_6_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2744_nl = MUX_s_1_2_2(buf_acc_data_11_13_0_sva,
      buf_acc_data_11_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2744_nl,
      buf_acc_data_11_13_0_sva, or_dcpl_124);
  assign buf_acc_data_11_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_13_45_1_sva_dfm_1,
      buf_acc_data_11_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_13_56_46_sva_dfm_1,
      buf_acc_data_11_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2746_nl = MUX_s_1_2_2(buf_acc_data_6_4_0_sva,
      buf_acc_data_6_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2746_nl,
      buf_acc_data_6_4_0_sva, or_dcpl_124);
  assign buf_acc_data_6_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_4_45_1_sva_dfm_1,
      buf_acc_data_6_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_4_56_46_sva_dfm_1,
      buf_acc_data_6_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2748_nl = MUX_s_1_2_2(buf_acc_data_11_12_0_sva,
      buf_acc_data_11_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2748_nl,
      buf_acc_data_11_12_0_sva, or_dcpl_124);
  assign buf_acc_data_11_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_12_45_1_sva_dfm_1,
      buf_acc_data_11_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_12_56_46_sva_dfm_1,
      buf_acc_data_11_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2750_nl = MUX_s_1_2_2(buf_acc_data_6_5_0_sva,
      buf_acc_data_6_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2750_nl,
      buf_acc_data_6_5_0_sva, or_dcpl_124);
  assign buf_acc_data_6_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_5_45_1_sva_dfm_1,
      buf_acc_data_6_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_5_56_46_sva_dfm_1,
      buf_acc_data_6_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2752_nl = MUX_s_1_2_2(buf_acc_data_11_11_0_sva,
      buf_acc_data_11_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2752_nl,
      buf_acc_data_11_11_0_sva, or_dcpl_124);
  assign buf_acc_data_11_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_11_45_1_sva_dfm_1,
      buf_acc_data_11_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_11_56_46_sva_dfm_1,
      buf_acc_data_11_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2754_nl = MUX_s_1_2_2(buf_acc_data_6_6_0_sva,
      buf_acc_data_6_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2754_nl,
      buf_acc_data_6_6_0_sva, or_dcpl_124);
  assign buf_acc_data_6_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_6_45_1_sva_dfm_1,
      buf_acc_data_6_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_6_56_46_sva_dfm_1,
      buf_acc_data_6_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2756_nl = MUX_s_1_2_2(buf_acc_data_11_10_0_sva,
      buf_acc_data_11_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2756_nl,
      buf_acc_data_11_10_0_sva, or_dcpl_124);
  assign buf_acc_data_11_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_10_45_1_sva_dfm_1,
      buf_acc_data_11_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_10_56_46_sva_dfm_1,
      buf_acc_data_11_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2758_nl = MUX_s_1_2_2(buf_acc_data_6_7_0_sva,
      buf_acc_data_6_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2758_nl,
      buf_acc_data_6_7_0_sva, or_dcpl_124);
  assign buf_acc_data_6_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_7_45_1_sva_dfm_1,
      buf_acc_data_6_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_7_56_46_sva_dfm_1,
      buf_acc_data_6_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2760_nl = MUX_s_1_2_2(buf_acc_data_11_9_0_sva,
      buf_acc_data_11_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2760_nl,
      buf_acc_data_11_9_0_sva, or_dcpl_124);
  assign buf_acc_data_11_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_9_45_1_sva_dfm_1,
      buf_acc_data_11_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_9_56_46_sva_dfm_1,
      buf_acc_data_11_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2762_nl = MUX_s_1_2_2(buf_acc_data_6_8_0_sva,
      buf_acc_data_6_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2762_nl,
      buf_acc_data_6_8_0_sva, or_dcpl_124);
  assign buf_acc_data_6_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_8_45_1_sva_dfm_1,
      buf_acc_data_6_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_8_56_46_sva_dfm_1,
      buf_acc_data_6_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2764_nl = MUX_s_1_2_2(buf_acc_data_11_8_0_sva,
      buf_acc_data_11_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2764_nl,
      buf_acc_data_11_8_0_sva, or_dcpl_124);
  assign buf_acc_data_11_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_8_45_1_sva_dfm_1,
      buf_acc_data_11_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_8_56_46_sva_dfm_1,
      buf_acc_data_11_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2766_nl = MUX_s_1_2_2(buf_acc_data_6_9_0_sva,
      buf_acc_data_6_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2766_nl,
      buf_acc_data_6_9_0_sva, or_dcpl_124);
  assign buf_acc_data_6_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_9_45_1_sva_dfm_1,
      buf_acc_data_6_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_9_56_46_sva_dfm_1,
      buf_acc_data_6_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2768_nl = MUX_s_1_2_2(buf_acc_data_11_7_0_sva,
      buf_acc_data_11_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2768_nl,
      buf_acc_data_11_7_0_sva, or_dcpl_124);
  assign buf_acc_data_11_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_7_45_1_sva_dfm_1,
      buf_acc_data_11_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_7_56_46_sva_dfm_1,
      buf_acc_data_11_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2770_nl = MUX_s_1_2_2(buf_acc_data_6_10_0_sva,
      buf_acc_data_6_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2770_nl,
      buf_acc_data_6_10_0_sva, or_dcpl_124);
  assign buf_acc_data_6_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_10_45_1_sva_dfm_1,
      buf_acc_data_6_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_10_56_46_sva_dfm_1,
      buf_acc_data_6_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2772_nl = MUX_s_1_2_2(buf_acc_data_11_6_0_sva,
      buf_acc_data_11_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2772_nl,
      buf_acc_data_11_6_0_sva, or_dcpl_124);
  assign buf_acc_data_11_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_6_45_1_sva_dfm_1,
      buf_acc_data_11_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_6_56_46_sva_dfm_1,
      buf_acc_data_11_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2774_nl = MUX_s_1_2_2(buf_acc_data_6_11_0_sva,
      buf_acc_data_6_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2774_nl,
      buf_acc_data_6_11_0_sva, or_dcpl_124);
  assign buf_acc_data_6_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_11_45_1_sva_dfm_1,
      buf_acc_data_6_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_11_56_46_sva_dfm_1,
      buf_acc_data_6_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2776_nl = MUX_s_1_2_2(buf_acc_data_11_5_0_sva,
      buf_acc_data_11_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2776_nl,
      buf_acc_data_11_5_0_sva, or_dcpl_124);
  assign buf_acc_data_11_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_5_45_1_sva_dfm_1,
      buf_acc_data_11_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_5_56_46_sva_dfm_1,
      buf_acc_data_11_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2778_nl = MUX_s_1_2_2(buf_acc_data_6_12_0_sva,
      buf_acc_data_6_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2778_nl,
      buf_acc_data_6_12_0_sva, or_dcpl_124);
  assign buf_acc_data_6_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_12_45_1_sva_dfm_1,
      buf_acc_data_6_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_12_56_46_sva_dfm_1,
      buf_acc_data_6_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2780_nl = MUX_s_1_2_2(buf_acc_data_11_4_0_sva,
      buf_acc_data_11_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2780_nl,
      buf_acc_data_11_4_0_sva, or_dcpl_124);
  assign buf_acc_data_11_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_4_45_1_sva_dfm_1,
      buf_acc_data_11_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_4_56_46_sva_dfm_1,
      buf_acc_data_11_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2782_nl = MUX_s_1_2_2(buf_acc_data_6_13_0_sva,
      buf_acc_data_6_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2782_nl,
      buf_acc_data_6_13_0_sva, or_dcpl_124);
  assign buf_acc_data_6_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_13_45_1_sva_dfm_1,
      buf_acc_data_6_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_13_56_46_sva_dfm_1,
      buf_acc_data_6_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2784_nl = MUX_s_1_2_2(buf_acc_data_11_3_0_sva,
      buf_acc_data_11_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2784_nl,
      buf_acc_data_11_3_0_sva, or_dcpl_124);
  assign buf_acc_data_11_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_3_45_1_sva_dfm_1,
      buf_acc_data_11_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_3_56_46_sva_dfm_1,
      buf_acc_data_11_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2786_nl = MUX_s_1_2_2(buf_acc_data_6_14_0_sva,
      buf_acc_data_6_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2786_nl,
      buf_acc_data_6_14_0_sva, or_dcpl_124);
  assign buf_acc_data_6_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_14_45_1_sva_dfm_1,
      buf_acc_data_6_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_14_56_46_sva_dfm_1,
      buf_acc_data_6_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2788_nl = MUX_s_1_2_2(buf_acc_data_11_2_0_sva,
      buf_acc_data_11_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2788_nl,
      buf_acc_data_11_2_0_sva, or_dcpl_124);
  assign buf_acc_data_11_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_2_45_1_sva_dfm_1,
      buf_acc_data_11_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_2_56_46_sva_dfm_1,
      buf_acc_data_11_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2790_nl = MUX_s_1_2_2(buf_acc_data_6_15_0_sva,
      buf_acc_data_6_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2790_nl,
      buf_acc_data_6_15_0_sva, or_dcpl_124);
  assign buf_acc_data_6_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_15_45_1_sva_dfm_1,
      buf_acc_data_6_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_15_56_46_sva_dfm_1,
      buf_acc_data_6_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2792_nl = MUX_s_1_2_2(buf_acc_data_11_1_0_sva,
      buf_acc_data_11_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2792_nl,
      buf_acc_data_11_1_0_sva, or_dcpl_124);
  assign buf_acc_data_11_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_1_45_1_sva_dfm_1,
      buf_acc_data_11_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_1_56_46_sva_dfm_1,
      buf_acc_data_11_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2794_nl = MUX_s_1_2_2(buf_acc_data_6_16_0_sva,
      buf_acc_data_6_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2794_nl,
      buf_acc_data_6_16_0_sva, or_dcpl_124);
  assign buf_acc_data_6_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_16_45_1_sva_dfm_1,
      buf_acc_data_6_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_16_56_46_sva_dfm_1,
      buf_acc_data_6_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2796_nl = MUX_s_1_2_2(buf_acc_data_11_0_0_sva,
      buf_acc_data_11_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_11_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2796_nl,
      buf_acc_data_11_0_0_sva, or_dcpl_124);
  assign buf_acc_data_11_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_11_0_45_1_sva_dfm_1,
      buf_acc_data_11_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_11_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_11_0_56_46_sva_dfm_1,
      buf_acc_data_11_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2798_nl = MUX_s_1_2_2(buf_acc_data_6_17_0_sva,
      buf_acc_data_6_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_6_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2798_nl,
      buf_acc_data_6_17_0_sva, or_dcpl_124);
  assign buf_acc_data_6_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_6_17_45_1_sva_dfm_1,
      buf_acc_data_6_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_6_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_6_17_56_46_sva_dfm_1,
      buf_acc_data_6_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2800_nl = MUX_s_1_2_2(buf_acc_data_10_17_0_sva,
      buf_acc_data_10_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2800_nl,
      buf_acc_data_10_17_0_sva, or_dcpl_124);
  assign buf_acc_data_10_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_17_45_1_sva_dfm_1,
      buf_acc_data_10_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_17_56_46_sva_dfm_1,
      buf_acc_data_10_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2802_nl = MUX_s_1_2_2(buf_acc_data_7_0_0_sva,
      buf_acc_data_7_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2802_nl,
      buf_acc_data_7_0_0_sva, or_dcpl_124);
  assign buf_acc_data_7_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_0_45_1_sva_dfm_1,
      buf_acc_data_7_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_0_56_46_sva_dfm_1,
      buf_acc_data_7_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2804_nl = MUX_s_1_2_2(buf_acc_data_10_16_0_sva,
      buf_acc_data_10_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2804_nl,
      buf_acc_data_10_16_0_sva, or_dcpl_124);
  assign buf_acc_data_10_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_16_45_1_sva_dfm_1,
      buf_acc_data_10_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_16_56_46_sva_dfm_1,
      buf_acc_data_10_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2806_nl = MUX_s_1_2_2(buf_acc_data_7_1_0_sva,
      buf_acc_data_7_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2806_nl,
      buf_acc_data_7_1_0_sva, or_dcpl_124);
  assign buf_acc_data_7_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_1_45_1_sva_dfm_1,
      buf_acc_data_7_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_1_56_46_sva_dfm_1,
      buf_acc_data_7_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2808_nl = MUX_s_1_2_2(buf_acc_data_10_15_0_sva,
      buf_acc_data_10_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2808_nl,
      buf_acc_data_10_15_0_sva, or_dcpl_124);
  assign buf_acc_data_10_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_15_45_1_sva_dfm_1,
      buf_acc_data_10_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_15_56_46_sva_dfm_1,
      buf_acc_data_10_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2810_nl = MUX_s_1_2_2(buf_acc_data_7_2_0_sva,
      buf_acc_data_7_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2810_nl,
      buf_acc_data_7_2_0_sva, or_dcpl_124);
  assign buf_acc_data_7_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_2_45_1_sva_dfm_1,
      buf_acc_data_7_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_2_56_46_sva_dfm_1,
      buf_acc_data_7_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2812_nl = MUX_s_1_2_2(buf_acc_data_10_14_0_sva,
      buf_acc_data_10_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2812_nl,
      buf_acc_data_10_14_0_sva, or_dcpl_124);
  assign buf_acc_data_10_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_14_45_1_sva_dfm_1,
      buf_acc_data_10_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_14_56_46_sva_dfm_1,
      buf_acc_data_10_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2814_nl = MUX_s_1_2_2(buf_acc_data_7_3_0_sva,
      buf_acc_data_7_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2814_nl,
      buf_acc_data_7_3_0_sva, or_dcpl_124);
  assign buf_acc_data_7_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_3_45_1_sva_dfm_1,
      buf_acc_data_7_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_3_56_46_sva_dfm_1,
      buf_acc_data_7_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2816_nl = MUX_s_1_2_2(buf_acc_data_10_13_0_sva,
      buf_acc_data_10_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2816_nl,
      buf_acc_data_10_13_0_sva, or_dcpl_124);
  assign buf_acc_data_10_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_13_45_1_sva_dfm_1,
      buf_acc_data_10_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_13_56_46_sva_dfm_1,
      buf_acc_data_10_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2818_nl = MUX_s_1_2_2(buf_acc_data_7_4_0_sva,
      buf_acc_data_7_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2818_nl,
      buf_acc_data_7_4_0_sva, or_dcpl_124);
  assign buf_acc_data_7_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_4_45_1_sva_dfm_1,
      buf_acc_data_7_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_4_56_46_sva_dfm_1,
      buf_acc_data_7_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2820_nl = MUX_s_1_2_2(buf_acc_data_10_12_0_sva,
      buf_acc_data_10_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2820_nl,
      buf_acc_data_10_12_0_sva, or_dcpl_124);
  assign buf_acc_data_10_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_12_45_1_sva_dfm_1,
      buf_acc_data_10_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_12_56_46_sva_dfm_1,
      buf_acc_data_10_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2822_nl = MUX_s_1_2_2(buf_acc_data_7_5_0_sva,
      buf_acc_data_7_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2822_nl,
      buf_acc_data_7_5_0_sva, or_dcpl_124);
  assign buf_acc_data_7_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_5_45_1_sva_dfm_1,
      buf_acc_data_7_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_5_56_46_sva_dfm_1,
      buf_acc_data_7_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2824_nl = MUX_s_1_2_2(buf_acc_data_10_11_0_sva,
      buf_acc_data_10_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2824_nl,
      buf_acc_data_10_11_0_sva, or_dcpl_124);
  assign buf_acc_data_10_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_11_45_1_sva_dfm_1,
      buf_acc_data_10_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_11_56_46_sva_dfm_1,
      buf_acc_data_10_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2826_nl = MUX_s_1_2_2(buf_acc_data_7_6_0_sva,
      buf_acc_data_7_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2826_nl,
      buf_acc_data_7_6_0_sva, or_dcpl_124);
  assign buf_acc_data_7_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_6_45_1_sva_dfm_1,
      buf_acc_data_7_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_6_56_46_sva_dfm_1,
      buf_acc_data_7_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2828_nl = MUX_s_1_2_2(buf_acc_data_10_10_0_sva,
      buf_acc_data_10_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2828_nl,
      buf_acc_data_10_10_0_sva, or_dcpl_124);
  assign buf_acc_data_10_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_10_45_1_sva_dfm_1,
      buf_acc_data_10_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_10_56_46_sva_dfm_1,
      buf_acc_data_10_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2830_nl = MUX_s_1_2_2(buf_acc_data_7_7_0_sva,
      buf_acc_data_7_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2830_nl,
      buf_acc_data_7_7_0_sva, or_dcpl_124);
  assign buf_acc_data_7_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_7_45_1_sva_dfm_1,
      buf_acc_data_7_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_7_56_46_sva_dfm_1,
      buf_acc_data_7_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2832_nl = MUX_s_1_2_2(buf_acc_data_10_9_0_sva,
      buf_acc_data_10_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2832_nl,
      buf_acc_data_10_9_0_sva, or_dcpl_124);
  assign buf_acc_data_10_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_9_45_1_sva_dfm_1,
      buf_acc_data_10_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_9_56_46_sva_dfm_1,
      buf_acc_data_10_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2834_nl = MUX_s_1_2_2(buf_acc_data_7_8_0_sva,
      buf_acc_data_7_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2834_nl,
      buf_acc_data_7_8_0_sva, or_dcpl_124);
  assign buf_acc_data_7_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_8_45_1_sva_dfm_1,
      buf_acc_data_7_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_8_56_46_sva_dfm_1,
      buf_acc_data_7_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2836_nl = MUX_s_1_2_2(buf_acc_data_10_8_0_sva,
      buf_acc_data_10_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2836_nl,
      buf_acc_data_10_8_0_sva, or_dcpl_124);
  assign buf_acc_data_10_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_8_45_1_sva_dfm_1,
      buf_acc_data_10_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_8_56_46_sva_dfm_1,
      buf_acc_data_10_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2838_nl = MUX_s_1_2_2(buf_acc_data_7_9_0_sva,
      buf_acc_data_7_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2838_nl,
      buf_acc_data_7_9_0_sva, or_dcpl_124);
  assign buf_acc_data_7_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_9_45_1_sva_dfm_1,
      buf_acc_data_7_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_9_56_46_sva_dfm_1,
      buf_acc_data_7_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2840_nl = MUX_s_1_2_2(buf_acc_data_10_7_0_sva,
      buf_acc_data_10_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2840_nl,
      buf_acc_data_10_7_0_sva, or_dcpl_124);
  assign buf_acc_data_10_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_7_45_1_sva_dfm_1,
      buf_acc_data_10_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_7_56_46_sva_dfm_1,
      buf_acc_data_10_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2842_nl = MUX_s_1_2_2(buf_acc_data_7_10_0_sva,
      buf_acc_data_7_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2842_nl,
      buf_acc_data_7_10_0_sva, or_dcpl_124);
  assign buf_acc_data_7_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_10_45_1_sva_dfm_1,
      buf_acc_data_7_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_10_56_46_sva_dfm_1,
      buf_acc_data_7_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2844_nl = MUX_s_1_2_2(buf_acc_data_10_6_0_sva,
      buf_acc_data_10_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2844_nl,
      buf_acc_data_10_6_0_sva, or_dcpl_124);
  assign buf_acc_data_10_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_6_45_1_sva_dfm_1,
      buf_acc_data_10_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_6_56_46_sva_dfm_1,
      buf_acc_data_10_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2846_nl = MUX_s_1_2_2(buf_acc_data_7_11_0_sva,
      buf_acc_data_7_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2846_nl,
      buf_acc_data_7_11_0_sva, or_dcpl_124);
  assign buf_acc_data_7_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_11_45_1_sva_dfm_1,
      buf_acc_data_7_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_11_56_46_sva_dfm_1,
      buf_acc_data_7_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2848_nl = MUX_s_1_2_2(buf_acc_data_10_5_0_sva,
      buf_acc_data_10_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2848_nl,
      buf_acc_data_10_5_0_sva, or_dcpl_124);
  assign buf_acc_data_10_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_5_45_1_sva_dfm_1,
      buf_acc_data_10_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_5_56_46_sva_dfm_1,
      buf_acc_data_10_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2850_nl = MUX_s_1_2_2(buf_acc_data_7_12_0_sva,
      buf_acc_data_7_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2850_nl,
      buf_acc_data_7_12_0_sva, or_dcpl_124);
  assign buf_acc_data_7_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_12_45_1_sva_dfm_1,
      buf_acc_data_7_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_12_56_46_sva_dfm_1,
      buf_acc_data_7_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2852_nl = MUX_s_1_2_2(buf_acc_data_10_4_0_sva,
      buf_acc_data_10_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2852_nl,
      buf_acc_data_10_4_0_sva, or_dcpl_124);
  assign buf_acc_data_10_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_4_45_1_sva_dfm_1,
      buf_acc_data_10_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_4_56_46_sva_dfm_1,
      buf_acc_data_10_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2854_nl = MUX_s_1_2_2(buf_acc_data_7_13_0_sva,
      buf_acc_data_7_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2854_nl,
      buf_acc_data_7_13_0_sva, or_dcpl_124);
  assign buf_acc_data_7_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_13_45_1_sva_dfm_1,
      buf_acc_data_7_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_13_56_46_sva_dfm_1,
      buf_acc_data_7_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2856_nl = MUX_s_1_2_2(buf_acc_data_10_3_0_sva,
      buf_acc_data_10_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2856_nl,
      buf_acc_data_10_3_0_sva, or_dcpl_124);
  assign buf_acc_data_10_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_3_45_1_sva_dfm_1,
      buf_acc_data_10_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_3_56_46_sva_dfm_1,
      buf_acc_data_10_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2858_nl = MUX_s_1_2_2(buf_acc_data_7_14_0_sva,
      buf_acc_data_7_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2858_nl,
      buf_acc_data_7_14_0_sva, or_dcpl_124);
  assign buf_acc_data_7_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_14_45_1_sva_dfm_1,
      buf_acc_data_7_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_14_56_46_sva_dfm_1,
      buf_acc_data_7_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2860_nl = MUX_s_1_2_2(buf_acc_data_10_2_0_sva,
      buf_acc_data_10_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2860_nl,
      buf_acc_data_10_2_0_sva, or_dcpl_124);
  assign buf_acc_data_10_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_2_45_1_sva_dfm_1,
      buf_acc_data_10_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_2_56_46_sva_dfm_1,
      buf_acc_data_10_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2862_nl = MUX_s_1_2_2(buf_acc_data_7_15_0_sva,
      buf_acc_data_7_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2862_nl,
      buf_acc_data_7_15_0_sva, or_dcpl_124);
  assign buf_acc_data_7_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_15_45_1_sva_dfm_1,
      buf_acc_data_7_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_15_56_46_sva_dfm_1,
      buf_acc_data_7_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2864_nl = MUX_s_1_2_2(buf_acc_data_10_1_0_sva,
      buf_acc_data_10_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2864_nl,
      buf_acc_data_10_1_0_sva, or_dcpl_124);
  assign buf_acc_data_10_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_1_45_1_sva_dfm_1,
      buf_acc_data_10_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_1_56_46_sva_dfm_1,
      buf_acc_data_10_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2866_nl = MUX_s_1_2_2(buf_acc_data_7_16_0_sva,
      buf_acc_data_7_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2866_nl,
      buf_acc_data_7_16_0_sva, or_dcpl_124);
  assign buf_acc_data_7_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_16_45_1_sva_dfm_1,
      buf_acc_data_7_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_16_56_46_sva_dfm_1,
      buf_acc_data_7_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2868_nl = MUX_s_1_2_2(buf_acc_data_10_0_0_sva,
      buf_acc_data_10_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_10_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2868_nl,
      buf_acc_data_10_0_0_sva, or_dcpl_124);
  assign buf_acc_data_10_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_10_0_45_1_sva_dfm_1,
      buf_acc_data_10_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_10_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_10_0_56_46_sva_dfm_1,
      buf_acc_data_10_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2870_nl = MUX_s_1_2_2(buf_acc_data_7_17_0_sva,
      buf_acc_data_7_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_7_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2870_nl,
      buf_acc_data_7_17_0_sva, or_dcpl_124);
  assign buf_acc_data_7_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_7_17_45_1_sva_dfm_1,
      buf_acc_data_7_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_7_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_7_17_56_46_sva_dfm_1,
      buf_acc_data_7_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2872_nl = MUX_s_1_2_2(buf_acc_data_9_17_0_sva,
      buf_acc_data_9_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2872_nl,
      buf_acc_data_9_17_0_sva, or_dcpl_124);
  assign buf_acc_data_9_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_17_45_1_sva_dfm_1,
      buf_acc_data_9_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_17_56_46_sva_dfm_1,
      buf_acc_data_9_17_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2874_nl = MUX_s_1_2_2(buf_acc_data_8_0_0_sva,
      buf_acc_data_8_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2874_nl,
      buf_acc_data_8_0_0_sva, or_dcpl_124);
  assign buf_acc_data_8_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_0_45_1_sva_dfm_1,
      buf_acc_data_8_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_0_56_46_sva_dfm_1,
      buf_acc_data_8_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2876_nl = MUX_s_1_2_2(buf_acc_data_9_16_0_sva,
      buf_acc_data_9_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2876_nl,
      buf_acc_data_9_16_0_sva, or_dcpl_124);
  assign buf_acc_data_9_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_16_45_1_sva_dfm_1,
      buf_acc_data_9_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_16_56_46_sva_dfm_1,
      buf_acc_data_9_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2878_nl = MUX_s_1_2_2(buf_acc_data_8_1_0_sva,
      buf_acc_data_8_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2878_nl,
      buf_acc_data_8_1_0_sva, or_dcpl_124);
  assign buf_acc_data_8_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_1_45_1_sva_dfm_1,
      buf_acc_data_8_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_1_56_46_sva_dfm_1,
      buf_acc_data_8_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2880_nl = MUX_s_1_2_2(buf_acc_data_9_15_0_sva,
      buf_acc_data_9_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2880_nl,
      buf_acc_data_9_15_0_sva, or_dcpl_124);
  assign buf_acc_data_9_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_15_45_1_sva_dfm_1,
      buf_acc_data_9_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_15_56_46_sva_dfm_1,
      buf_acc_data_9_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2882_nl = MUX_s_1_2_2(buf_acc_data_8_2_0_sva,
      buf_acc_data_8_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2882_nl,
      buf_acc_data_8_2_0_sva, or_dcpl_124);
  assign buf_acc_data_8_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_2_45_1_sva_dfm_1,
      buf_acc_data_8_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_2_56_46_sva_dfm_1,
      buf_acc_data_8_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2884_nl = MUX_s_1_2_2(buf_acc_data_9_14_0_sva,
      buf_acc_data_9_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2884_nl,
      buf_acc_data_9_14_0_sva, or_dcpl_124);
  assign buf_acc_data_9_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_14_45_1_sva_dfm_1,
      buf_acc_data_9_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_14_56_46_sva_dfm_1,
      buf_acc_data_9_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2886_nl = MUX_s_1_2_2(buf_acc_data_8_3_0_sva,
      buf_acc_data_8_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2886_nl,
      buf_acc_data_8_3_0_sva, or_dcpl_124);
  assign buf_acc_data_8_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_3_45_1_sva_dfm_1,
      buf_acc_data_8_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_3_56_46_sva_dfm_1,
      buf_acc_data_8_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2888_nl = MUX_s_1_2_2(buf_acc_data_9_13_0_sva,
      buf_acc_data_9_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2888_nl,
      buf_acc_data_9_13_0_sva, or_dcpl_124);
  assign buf_acc_data_9_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_13_45_1_sva_dfm_1,
      buf_acc_data_9_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_13_56_46_sva_dfm_1,
      buf_acc_data_9_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2890_nl = MUX_s_1_2_2(buf_acc_data_8_4_0_sva,
      buf_acc_data_8_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2890_nl,
      buf_acc_data_8_4_0_sva, or_dcpl_124);
  assign buf_acc_data_8_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_4_45_1_sva_dfm_1,
      buf_acc_data_8_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_4_56_46_sva_dfm_1,
      buf_acc_data_8_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2892_nl = MUX_s_1_2_2(buf_acc_data_9_12_0_sva,
      buf_acc_data_9_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2892_nl,
      buf_acc_data_9_12_0_sva, or_dcpl_124);
  assign buf_acc_data_9_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_12_45_1_sva_dfm_1,
      buf_acc_data_9_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_12_56_46_sva_dfm_1,
      buf_acc_data_9_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2894_nl = MUX_s_1_2_2(buf_acc_data_8_5_0_sva,
      buf_acc_data_8_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2894_nl,
      buf_acc_data_8_5_0_sva, or_dcpl_124);
  assign buf_acc_data_8_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_5_45_1_sva_dfm_1,
      buf_acc_data_8_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_5_56_46_sva_dfm_1,
      buf_acc_data_8_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2896_nl = MUX_s_1_2_2(buf_acc_data_9_11_0_sva,
      buf_acc_data_9_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2896_nl,
      buf_acc_data_9_11_0_sva, or_dcpl_124);
  assign buf_acc_data_9_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_11_45_1_sva_dfm_1,
      buf_acc_data_9_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_11_56_46_sva_dfm_1,
      buf_acc_data_9_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2898_nl = MUX_s_1_2_2(buf_acc_data_8_6_0_sva,
      buf_acc_data_8_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2898_nl,
      buf_acc_data_8_6_0_sva, or_dcpl_124);
  assign buf_acc_data_8_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_6_45_1_sva_dfm_1,
      buf_acc_data_8_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_6_56_46_sva_dfm_1,
      buf_acc_data_8_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2900_nl = MUX_s_1_2_2(buf_acc_data_9_10_0_sva,
      buf_acc_data_9_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2900_nl,
      buf_acc_data_9_10_0_sva, or_dcpl_124);
  assign buf_acc_data_9_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_10_45_1_sva_dfm_1,
      buf_acc_data_9_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_10_56_46_sva_dfm_1,
      buf_acc_data_9_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2902_nl = MUX_s_1_2_2(buf_acc_data_8_7_0_sva,
      buf_acc_data_8_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2902_nl,
      buf_acc_data_8_7_0_sva, or_dcpl_124);
  assign buf_acc_data_8_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_7_45_1_sva_dfm_1,
      buf_acc_data_8_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_7_56_46_sva_dfm_1,
      buf_acc_data_8_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2904_nl = MUX_s_1_2_2(buf_acc_data_9_9_0_sva,
      buf_acc_data_9_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2904_nl,
      buf_acc_data_9_9_0_sva, or_dcpl_124);
  assign buf_acc_data_9_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_9_45_1_sva_dfm_1,
      buf_acc_data_9_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_9_56_46_sva_dfm_1,
      buf_acc_data_9_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2906_nl = MUX_s_1_2_2(buf_acc_data_8_8_0_sva,
      buf_acc_data_8_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2906_nl,
      buf_acc_data_8_8_0_sva, or_dcpl_124);
  assign buf_acc_data_8_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_8_45_1_sva_dfm_1,
      buf_acc_data_8_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_8_56_46_sva_dfm_1,
      buf_acc_data_8_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2908_nl = MUX_s_1_2_2(buf_acc_data_9_8_0_sva,
      buf_acc_data_9_8_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_8_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2908_nl,
      buf_acc_data_9_8_0_sva, or_dcpl_124);
  assign buf_acc_data_9_8_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_8_45_1_sva_dfm_1,
      buf_acc_data_9_8_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_8_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_8_56_46_sva_dfm_1,
      buf_acc_data_9_8_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2910_nl = MUX_s_1_2_2(buf_acc_data_8_9_0_sva,
      buf_acc_data_8_9_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_9_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2910_nl,
      buf_acc_data_8_9_0_sva, or_dcpl_124);
  assign buf_acc_data_8_9_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_9_45_1_sva_dfm_1,
      buf_acc_data_8_9_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_9_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_9_56_46_sva_dfm_1,
      buf_acc_data_8_9_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2912_nl = MUX_s_1_2_2(buf_acc_data_9_7_0_sva,
      buf_acc_data_9_7_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_7_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2912_nl,
      buf_acc_data_9_7_0_sva, or_dcpl_124);
  assign buf_acc_data_9_7_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_7_45_1_sva_dfm_1,
      buf_acc_data_9_7_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_7_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_7_56_46_sva_dfm_1,
      buf_acc_data_9_7_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2914_nl = MUX_s_1_2_2(buf_acc_data_8_10_0_sva,
      buf_acc_data_8_10_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_10_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2914_nl,
      buf_acc_data_8_10_0_sva, or_dcpl_124);
  assign buf_acc_data_8_10_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_10_45_1_sva_dfm_1,
      buf_acc_data_8_10_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_10_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_10_56_46_sva_dfm_1,
      buf_acc_data_8_10_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2916_nl = MUX_s_1_2_2(buf_acc_data_9_6_0_sva,
      buf_acc_data_9_6_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_6_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2916_nl,
      buf_acc_data_9_6_0_sva, or_dcpl_124);
  assign buf_acc_data_9_6_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_6_45_1_sva_dfm_1,
      buf_acc_data_9_6_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_6_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_6_56_46_sva_dfm_1,
      buf_acc_data_9_6_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2918_nl = MUX_s_1_2_2(buf_acc_data_8_11_0_sva,
      buf_acc_data_8_11_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_11_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2918_nl,
      buf_acc_data_8_11_0_sva, or_dcpl_124);
  assign buf_acc_data_8_11_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_11_45_1_sva_dfm_1,
      buf_acc_data_8_11_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_11_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_11_56_46_sva_dfm_1,
      buf_acc_data_8_11_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2920_nl = MUX_s_1_2_2(buf_acc_data_9_5_0_sva,
      buf_acc_data_9_5_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_5_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2920_nl,
      buf_acc_data_9_5_0_sva, or_dcpl_124);
  assign buf_acc_data_9_5_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_5_45_1_sva_dfm_1,
      buf_acc_data_9_5_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_5_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_5_56_46_sva_dfm_1,
      buf_acc_data_9_5_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2922_nl = MUX_s_1_2_2(buf_acc_data_8_12_0_sva,
      buf_acc_data_8_12_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_12_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2922_nl,
      buf_acc_data_8_12_0_sva, or_dcpl_124);
  assign buf_acc_data_8_12_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_12_45_1_sva_dfm_1,
      buf_acc_data_8_12_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_12_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_12_56_46_sva_dfm_1,
      buf_acc_data_8_12_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2924_nl = MUX_s_1_2_2(buf_acc_data_9_4_0_sva,
      buf_acc_data_9_4_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_4_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2924_nl,
      buf_acc_data_9_4_0_sva, or_dcpl_124);
  assign buf_acc_data_9_4_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_4_45_1_sva_dfm_1,
      buf_acc_data_9_4_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_4_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_4_56_46_sva_dfm_1,
      buf_acc_data_9_4_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2926_nl = MUX_s_1_2_2(buf_acc_data_8_13_0_sva,
      buf_acc_data_8_13_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_13_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2926_nl,
      buf_acc_data_8_13_0_sva, or_dcpl_124);
  assign buf_acc_data_8_13_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_13_45_1_sva_dfm_1,
      buf_acc_data_8_13_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_13_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_13_56_46_sva_dfm_1,
      buf_acc_data_8_13_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2928_nl = MUX_s_1_2_2(buf_acc_data_9_3_0_sva,
      buf_acc_data_9_3_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_3_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2928_nl,
      buf_acc_data_9_3_0_sva, or_dcpl_124);
  assign buf_acc_data_9_3_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_3_45_1_sva_dfm_1,
      buf_acc_data_9_3_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_3_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_3_56_46_sva_dfm_1,
      buf_acc_data_9_3_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2930_nl = MUX_s_1_2_2(buf_acc_data_8_14_0_sva,
      buf_acc_data_8_14_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_14_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2930_nl,
      buf_acc_data_8_14_0_sva, or_dcpl_124);
  assign buf_acc_data_8_14_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_14_45_1_sva_dfm_1,
      buf_acc_data_8_14_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_14_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_14_56_46_sva_dfm_1,
      buf_acc_data_8_14_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2932_nl = MUX_s_1_2_2(buf_acc_data_9_2_0_sva,
      buf_acc_data_9_2_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_2_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2932_nl,
      buf_acc_data_9_2_0_sva, or_dcpl_124);
  assign buf_acc_data_9_2_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_2_45_1_sva_dfm_1,
      buf_acc_data_9_2_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_2_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_2_56_46_sva_dfm_1,
      buf_acc_data_9_2_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2934_nl = MUX_s_1_2_2(buf_acc_data_8_15_0_sva,
      buf_acc_data_8_15_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_15_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2934_nl,
      buf_acc_data_8_15_0_sva, or_dcpl_124);
  assign buf_acc_data_8_15_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_15_45_1_sva_dfm_1,
      buf_acc_data_8_15_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_15_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_15_56_46_sva_dfm_1,
      buf_acc_data_8_15_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2936_nl = MUX_s_1_2_2(buf_acc_data_9_1_0_sva,
      buf_acc_data_9_1_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_1_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2936_nl,
      buf_acc_data_9_1_0_sva, or_dcpl_124);
  assign buf_acc_data_9_1_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_1_45_1_sva_dfm_1,
      buf_acc_data_9_1_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_1_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_1_56_46_sva_dfm_1,
      buf_acc_data_9_1_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2938_nl = MUX_s_1_2_2(buf_acc_data_8_16_0_sva,
      buf_acc_data_8_16_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_16_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2938_nl,
      buf_acc_data_8_16_0_sva, or_dcpl_124);
  assign buf_acc_data_8_16_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_16_45_1_sva_dfm_1,
      buf_acc_data_8_16_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_16_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_16_56_46_sva_dfm_1,
      buf_acc_data_8_16_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2940_nl = MUX_s_1_2_2(buf_acc_data_9_0_0_sva,
      buf_acc_data_9_0_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_9_0_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2940_nl,
      buf_acc_data_9_0_0_sva, or_dcpl_124);
  assign buf_acc_data_9_0_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_9_0_45_1_sva_dfm_1,
      buf_acc_data_9_0_45_1_sva, or_dcpl_127);
  assign buf_acc_data_9_0_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_9_0_56_46_sva_dfm_1,
      buf_acc_data_9_0_56_46_sva, or_dcpl_127);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2942_nl = MUX_s_1_2_2(buf_acc_data_8_17_0_sva,
      buf_acc_data_8_17_0_sva_dfm_mx0, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2);
  assign buf_acc_data_8_17_0_sva_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_for_mux_2942_nl,
      buf_acc_data_8_17_0_sva, or_dcpl_124);
  assign buf_acc_data_8_17_45_1_sva_mx0 = MUX_v_45_2_2(buf_acc_data_8_17_45_1_sva_dfm_1,
      buf_acc_data_8_17_45_1_sva, or_dcpl_127);
  assign buf_acc_data_8_17_56_46_sva_mx0 = MUX_v_11_2_2(buf_acc_data_8_17_56_46_sva_dfm_1,
      buf_acc_data_8_17_56_46_sva, or_dcpl_127);
  assign STORE_LOOP_mux_29_nl = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, STORE_LOOP_equal_tmp_2_2);
  assign CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_mx1 = MUX_s_1_2_2(STORE_LOOP_mux_29_nl,
      CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2, or_dcpl_88);
  assign STORE_LOOP_mux_30_nl = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2,
      CONVOLUTION_LOOP_for_for_for_acc_46_sva_2, STORE_LOOP_equal_tmp_2_2);
  assign CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_mx1 = MUX_s_1_2_2(STORE_LOOP_mux_30_nl,
      CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2, or_dcpl_88);
  assign CONVOLUTION_LOOP_for_for_for_acc_0_sva_2 = ~((~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[0])
      | CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl = ~(MUX_v_45_2_2((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[45:1]),
      45'b111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2 = ~(MUX_v_45_2_2(CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl,
      45'b111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_acc_46_sva_2 = ~((~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[46])
      | CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1 = ~((~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[0])
      | CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_nor_1_nl = ~(MUX_v_55_2_2((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[55:1]),
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0 = ~(MUX_v_55_2_2(CONVOLUTION_LOOP_for_for_for_else_nor_1_nl,
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1 = ~(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0
      | (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0
      & (~ (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1 = (~ CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0)
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0
      & (CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0[0]);
  assign nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1 = conv_s2s_57_58({CONVOLUTION_LOOP_for_for_for_else_mux_itm_1
      , CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1 , CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1})
      + conv_s2s_47_58({CONVOLUTION_LOOP_for_for_for_acc_46_sva_2 , CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2
      , CONVOLUTION_LOOP_for_for_for_acc_0_sva_2});
  assign CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:0];
  assign CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:56]==2'b10);
  assign CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:56]!=2'b01));
  assign CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_45_1_1
      = MUX_v_45_324_2(buf_acc_data_0_0_45_1_sva_dfm_1, buf_acc_data_0_1_45_1_sva_dfm_1,
      buf_acc_data_0_2_45_1_sva_dfm_1, buf_acc_data_0_3_45_1_sva_dfm_1, buf_acc_data_0_4_45_1_sva_dfm_1,
      buf_acc_data_0_5_45_1_sva_dfm_1, buf_acc_data_0_6_45_1_sva_dfm_1, buf_acc_data_0_7_45_1_sva_dfm_1,
      buf_acc_data_0_8_45_1_sva_dfm_1, buf_acc_data_0_9_45_1_sva_dfm_1, buf_acc_data_0_10_45_1_sva_dfm_1,
      buf_acc_data_0_11_45_1_sva_dfm_1, buf_acc_data_0_12_45_1_sva_dfm_1, buf_acc_data_0_13_45_1_sva_dfm_1,
      buf_acc_data_0_14_45_1_sva_dfm_1, buf_acc_data_0_15_45_1_sva_dfm_1, buf_acc_data_0_16_45_1_sva_dfm_1,
      buf_acc_data_0_17_45_1_sva_dfm_1, buf_acc_data_1_0_45_1_sva_dfm_1, buf_acc_data_1_1_45_1_sva_dfm_1,
      buf_acc_data_1_2_45_1_sva_dfm_1, buf_acc_data_1_3_45_1_sva_dfm_1, buf_acc_data_1_4_45_1_sva_dfm_1,
      buf_acc_data_1_5_45_1_sva_dfm_1, buf_acc_data_1_6_45_1_sva_dfm_1, buf_acc_data_1_7_45_1_sva_dfm_1,
      buf_acc_data_1_8_45_1_sva_dfm_1, buf_acc_data_1_9_45_1_sva_dfm_1, buf_acc_data_1_10_45_1_sva_dfm_1,
      buf_acc_data_1_11_45_1_sva_dfm_1, buf_acc_data_1_12_45_1_sva_dfm_1, buf_acc_data_1_13_45_1_sva_dfm_1,
      buf_acc_data_1_14_45_1_sva_dfm_1, buf_acc_data_1_15_45_1_sva_dfm_1, buf_acc_data_1_16_45_1_sva_dfm_1,
      buf_acc_data_1_17_45_1_sva_dfm_1, buf_acc_data_2_0_45_1_sva_dfm_1, buf_acc_data_2_1_45_1_sva_dfm_1,
      buf_acc_data_2_2_45_1_sva_dfm_1, buf_acc_data_2_3_45_1_sva_dfm_1, buf_acc_data_2_4_45_1_sva_dfm_1,
      buf_acc_data_2_5_45_1_sva_dfm_1, buf_acc_data_2_6_45_1_sva_dfm_1, buf_acc_data_2_7_45_1_sva_dfm_1,
      buf_acc_data_2_8_45_1_sva_dfm_1, buf_acc_data_2_9_45_1_sva_dfm_1, buf_acc_data_2_10_45_1_sva_dfm_1,
      buf_acc_data_2_11_45_1_sva_dfm_1, buf_acc_data_2_12_45_1_sva_dfm_1, buf_acc_data_2_13_45_1_sva_dfm_1,
      buf_acc_data_2_14_45_1_sva_dfm_1, buf_acc_data_2_15_45_1_sva_dfm_1, buf_acc_data_2_16_45_1_sva_dfm_1,
      buf_acc_data_2_17_45_1_sva_dfm_1, buf_acc_data_3_0_45_1_sva_dfm_1, buf_acc_data_3_1_45_1_sva_dfm_1,
      buf_acc_data_3_2_45_1_sva_dfm_1, buf_acc_data_3_3_45_1_sva_dfm_1, buf_acc_data_3_4_45_1_sva_dfm_1,
      buf_acc_data_3_5_45_1_sva_dfm_1, buf_acc_data_3_6_45_1_sva_dfm_1, buf_acc_data_3_7_45_1_sva_dfm_1,
      buf_acc_data_3_8_45_1_sva_dfm_1, buf_acc_data_3_9_45_1_sva_dfm_1, buf_acc_data_3_10_45_1_sva_dfm_1,
      buf_acc_data_3_11_45_1_sva_dfm_1, buf_acc_data_3_12_45_1_sva_dfm_1, buf_acc_data_3_13_45_1_sva_dfm_1,
      buf_acc_data_3_14_45_1_sva_dfm_1, buf_acc_data_3_15_45_1_sva_dfm_1, buf_acc_data_3_16_45_1_sva_dfm_1,
      buf_acc_data_3_17_45_1_sva_dfm_1, buf_acc_data_4_0_45_1_sva_dfm_1, buf_acc_data_4_1_45_1_sva_dfm_1,
      buf_acc_data_4_2_45_1_sva_dfm_1, buf_acc_data_4_3_45_1_sva_dfm_1, buf_acc_data_4_4_45_1_sva_dfm_1,
      buf_acc_data_4_5_45_1_sva_dfm_1, buf_acc_data_4_6_45_1_sva_dfm_1, buf_acc_data_4_7_45_1_sva_dfm_1,
      buf_acc_data_4_8_45_1_sva_dfm_1, buf_acc_data_4_9_45_1_sva_dfm_1, buf_acc_data_4_10_45_1_sva_dfm_1,
      buf_acc_data_4_11_45_1_sva_dfm_1, buf_acc_data_4_12_45_1_sva_dfm_1, buf_acc_data_4_13_45_1_sva_dfm_1,
      buf_acc_data_4_14_45_1_sva_dfm_1, buf_acc_data_4_15_45_1_sva_dfm_1, buf_acc_data_4_16_45_1_sva_dfm_1,
      buf_acc_data_4_17_45_1_sva_dfm_1, buf_acc_data_5_0_45_1_sva_dfm_1, buf_acc_data_5_1_45_1_sva_dfm_1,
      buf_acc_data_5_2_45_1_sva_dfm_1, buf_acc_data_5_3_45_1_sva_dfm_1, buf_acc_data_5_4_45_1_sva_dfm_1,
      buf_acc_data_5_5_45_1_sva_dfm_1, buf_acc_data_5_6_45_1_sva_dfm_1, buf_acc_data_5_7_45_1_sva_dfm_1,
      buf_acc_data_5_8_45_1_sva_dfm_1, buf_acc_data_5_9_45_1_sva_dfm_1, buf_acc_data_5_10_45_1_sva_dfm_1,
      buf_acc_data_5_11_45_1_sva_dfm_1, buf_acc_data_5_12_45_1_sva_dfm_1, buf_acc_data_5_13_45_1_sva_dfm_1,
      buf_acc_data_5_14_45_1_sva_dfm_1, buf_acc_data_5_15_45_1_sva_dfm_1, buf_acc_data_5_16_45_1_sva_dfm_1,
      buf_acc_data_5_17_45_1_sva_dfm_1, buf_acc_data_6_0_45_1_sva_dfm_1, buf_acc_data_6_1_45_1_sva_dfm_1,
      buf_acc_data_6_2_45_1_sva_dfm_1, buf_acc_data_6_3_45_1_sva_dfm_1, buf_acc_data_6_4_45_1_sva_dfm_1,
      buf_acc_data_6_5_45_1_sva_dfm_1, buf_acc_data_6_6_45_1_sva_dfm_1, buf_acc_data_6_7_45_1_sva_dfm_1,
      buf_acc_data_6_8_45_1_sva_dfm_1, buf_acc_data_6_9_45_1_sva_dfm_1, buf_acc_data_6_10_45_1_sva_dfm_1,
      buf_acc_data_6_11_45_1_sva_dfm_1, buf_acc_data_6_12_45_1_sva_dfm_1, buf_acc_data_6_13_45_1_sva_dfm_1,
      buf_acc_data_6_14_45_1_sva_dfm_1, buf_acc_data_6_15_45_1_sva_dfm_1, buf_acc_data_6_16_45_1_sva_dfm_1,
      buf_acc_data_6_17_45_1_sva_dfm_1, buf_acc_data_7_0_45_1_sva_dfm_1, buf_acc_data_7_1_45_1_sva_dfm_1,
      buf_acc_data_7_2_45_1_sva_dfm_1, buf_acc_data_7_3_45_1_sva_dfm_1, buf_acc_data_7_4_45_1_sva_dfm_1,
      buf_acc_data_7_5_45_1_sva_dfm_1, buf_acc_data_7_6_45_1_sva_dfm_1, buf_acc_data_7_7_45_1_sva_dfm_1,
      buf_acc_data_7_8_45_1_sva_dfm_1, buf_acc_data_7_9_45_1_sva_dfm_1, buf_acc_data_7_10_45_1_sva_dfm_1,
      buf_acc_data_7_11_45_1_sva_dfm_1, buf_acc_data_7_12_45_1_sva_dfm_1, buf_acc_data_7_13_45_1_sva_dfm_1,
      buf_acc_data_7_14_45_1_sva_dfm_1, buf_acc_data_7_15_45_1_sva_dfm_1, buf_acc_data_7_16_45_1_sva_dfm_1,
      buf_acc_data_7_17_45_1_sva_dfm_1, buf_acc_data_8_0_45_1_sva_dfm_1, buf_acc_data_8_1_45_1_sva_dfm_1,
      buf_acc_data_8_2_45_1_sva_dfm_1, buf_acc_data_8_3_45_1_sva_dfm_1, buf_acc_data_8_4_45_1_sva_dfm_1,
      buf_acc_data_8_5_45_1_sva_dfm_1, buf_acc_data_8_6_45_1_sva_dfm_1, buf_acc_data_8_7_45_1_sva_dfm_1,
      buf_acc_data_8_8_45_1_sva_dfm_1, buf_acc_data_8_9_45_1_sva_dfm_1, buf_acc_data_8_10_45_1_sva_dfm_1,
      buf_acc_data_8_11_45_1_sva_dfm_1, buf_acc_data_8_12_45_1_sva_dfm_1, buf_acc_data_8_13_45_1_sva_dfm_1,
      buf_acc_data_8_14_45_1_sva_dfm_1, buf_acc_data_8_15_45_1_sva_dfm_1, buf_acc_data_8_16_45_1_sva_dfm_1,
      buf_acc_data_8_17_45_1_sva_dfm_1, buf_acc_data_9_0_45_1_sva_dfm_1, buf_acc_data_9_1_45_1_sva_dfm_1,
      buf_acc_data_9_2_45_1_sva_dfm_1, buf_acc_data_9_3_45_1_sva_dfm_1, buf_acc_data_9_4_45_1_sva_dfm_1,
      buf_acc_data_9_5_45_1_sva_dfm_1, buf_acc_data_9_6_45_1_sva_dfm_1, buf_acc_data_9_7_45_1_sva_dfm_1,
      buf_acc_data_9_8_45_1_sva_dfm_1, buf_acc_data_9_9_45_1_sva_dfm_1, buf_acc_data_9_10_45_1_sva_dfm_1,
      buf_acc_data_9_11_45_1_sva_dfm_1, buf_acc_data_9_12_45_1_sva_dfm_1, buf_acc_data_9_13_45_1_sva_dfm_1,
      buf_acc_data_9_14_45_1_sva_dfm_1, buf_acc_data_9_15_45_1_sva_dfm_1, buf_acc_data_9_16_45_1_sva_dfm_1,
      buf_acc_data_9_17_45_1_sva_dfm_1, buf_acc_data_10_0_45_1_sva_dfm_1, buf_acc_data_10_1_45_1_sva_dfm_1,
      buf_acc_data_10_2_45_1_sva_dfm_1, buf_acc_data_10_3_45_1_sva_dfm_1, buf_acc_data_10_4_45_1_sva_dfm_1,
      buf_acc_data_10_5_45_1_sva_dfm_1, buf_acc_data_10_6_45_1_sva_dfm_1, buf_acc_data_10_7_45_1_sva_dfm_1,
      buf_acc_data_10_8_45_1_sva_dfm_1, buf_acc_data_10_9_45_1_sva_dfm_1, buf_acc_data_10_10_45_1_sva_dfm_1,
      buf_acc_data_10_11_45_1_sva_dfm_1, buf_acc_data_10_12_45_1_sva_dfm_1, buf_acc_data_10_13_45_1_sva_dfm_1,
      buf_acc_data_10_14_45_1_sva_dfm_1, buf_acc_data_10_15_45_1_sva_dfm_1, buf_acc_data_10_16_45_1_sva_dfm_1,
      buf_acc_data_10_17_45_1_sva_dfm_1, buf_acc_data_11_0_45_1_sva_dfm_1, buf_acc_data_11_1_45_1_sva_dfm_1,
      buf_acc_data_11_2_45_1_sva_dfm_1, buf_acc_data_11_3_45_1_sva_dfm_1, buf_acc_data_11_4_45_1_sva_dfm_1,
      buf_acc_data_11_5_45_1_sva_dfm_1, buf_acc_data_11_6_45_1_sva_dfm_1, buf_acc_data_11_7_45_1_sva_dfm_1,
      buf_acc_data_11_8_45_1_sva_dfm_1, buf_acc_data_11_9_45_1_sva_dfm_1, buf_acc_data_11_10_45_1_sva_dfm_1,
      buf_acc_data_11_11_45_1_sva_dfm_1, buf_acc_data_11_12_45_1_sva_dfm_1, buf_acc_data_11_13_45_1_sva_dfm_1,
      buf_acc_data_11_14_45_1_sva_dfm_1, buf_acc_data_11_15_45_1_sva_dfm_1, buf_acc_data_11_16_45_1_sva_dfm_1,
      buf_acc_data_11_17_45_1_sva_dfm_1, buf_acc_data_12_0_45_1_sva_dfm_1, buf_acc_data_12_1_45_1_sva_dfm_1,
      buf_acc_data_12_2_45_1_sva_dfm_1, buf_acc_data_12_3_45_1_sva_dfm_1, buf_acc_data_12_4_45_1_sva_dfm_1,
      buf_acc_data_12_5_45_1_sva_dfm_1, buf_acc_data_12_6_45_1_sva_dfm_1, buf_acc_data_12_7_45_1_sva_dfm_1,
      buf_acc_data_12_8_45_1_sva_dfm_1, buf_acc_data_12_9_45_1_sva_dfm_1, buf_acc_data_12_10_45_1_sva_dfm_1,
      buf_acc_data_12_11_45_1_sva_dfm_1, buf_acc_data_12_12_45_1_sva_dfm_1, buf_acc_data_12_13_45_1_sva_dfm_1,
      buf_acc_data_12_14_45_1_sva_dfm_1, buf_acc_data_12_15_45_1_sva_dfm_1, buf_acc_data_12_16_45_1_sva_dfm_1,
      buf_acc_data_12_17_45_1_sva_dfm_1, buf_acc_data_13_0_45_1_sva_dfm_1, buf_acc_data_13_1_45_1_sva_dfm_1,
      buf_acc_data_13_2_45_1_sva_dfm_1, buf_acc_data_13_3_45_1_sva_dfm_1, buf_acc_data_13_4_45_1_sva_dfm_1,
      buf_acc_data_13_5_45_1_sva_dfm_1, buf_acc_data_13_6_45_1_sva_dfm_1, buf_acc_data_13_7_45_1_sva_dfm_1,
      buf_acc_data_13_8_45_1_sva_dfm_1, buf_acc_data_13_9_45_1_sva_dfm_1, buf_acc_data_13_10_45_1_sva_dfm_1,
      buf_acc_data_13_11_45_1_sva_dfm_1, buf_acc_data_13_12_45_1_sva_dfm_1, buf_acc_data_13_13_45_1_sva_dfm_1,
      buf_acc_data_13_14_45_1_sva_dfm_1, buf_acc_data_13_15_45_1_sva_dfm_1, buf_acc_data_13_16_45_1_sva_dfm_1,
      buf_acc_data_13_17_45_1_sva_dfm_1, buf_acc_data_14_0_45_1_sva_dfm_1, buf_acc_data_14_1_45_1_sva_dfm_1,
      buf_acc_data_14_2_45_1_sva_dfm_1, buf_acc_data_14_3_45_1_sva_dfm_1, buf_acc_data_14_4_45_1_sva_dfm_1,
      buf_acc_data_14_5_45_1_sva_dfm_1, buf_acc_data_14_6_45_1_sva_dfm_1, buf_acc_data_14_7_45_1_sva_dfm_1,
      buf_acc_data_14_8_45_1_sva_dfm_1, buf_acc_data_14_9_45_1_sva_dfm_1, buf_acc_data_14_10_45_1_sva_dfm_1,
      buf_acc_data_14_11_45_1_sva_dfm_1, buf_acc_data_14_12_45_1_sva_dfm_1, buf_acc_data_14_13_45_1_sva_dfm_1,
      buf_acc_data_14_14_45_1_sva_dfm_1, buf_acc_data_14_15_45_1_sva_dfm_1, buf_acc_data_14_16_45_1_sva_dfm_1,
      buf_acc_data_14_17_45_1_sva_dfm_1, buf_acc_data_15_0_45_1_sva_dfm_1, buf_acc_data_15_1_45_1_sva_dfm_1,
      buf_acc_data_15_2_45_1_sva_dfm_1, buf_acc_data_15_3_45_1_sva_dfm_1, buf_acc_data_15_4_45_1_sva_dfm_1,
      buf_acc_data_15_5_45_1_sva_dfm_1, buf_acc_data_15_6_45_1_sva_dfm_1, buf_acc_data_15_7_45_1_sva_dfm_1,
      buf_acc_data_15_8_45_1_sva_dfm_1, buf_acc_data_15_9_45_1_sva_dfm_1, buf_acc_data_15_10_45_1_sva_dfm_1,
      buf_acc_data_15_11_45_1_sva_dfm_1, buf_acc_data_15_12_45_1_sva_dfm_1, buf_acc_data_15_13_45_1_sva_dfm_1,
      buf_acc_data_15_14_45_1_sva_dfm_1, buf_acc_data_15_15_45_1_sva_dfm_1, buf_acc_data_15_16_45_1_sva_dfm_1,
      buf_acc_data_15_17_45_1_sva_dfm_1, buf_acc_data_16_0_45_1_sva_dfm_1, buf_acc_data_16_1_45_1_sva_dfm_1,
      buf_acc_data_16_2_45_1_sva_dfm_1, buf_acc_data_16_3_45_1_sva_dfm_1, buf_acc_data_16_4_45_1_sva_dfm_1,
      buf_acc_data_16_5_45_1_sva_dfm_1, buf_acc_data_16_6_45_1_sva_dfm_1, buf_acc_data_16_7_45_1_sva_dfm_1,
      buf_acc_data_16_8_45_1_sva_dfm_1, buf_acc_data_16_9_45_1_sva_dfm_1, buf_acc_data_16_10_45_1_sva_dfm_1,
      buf_acc_data_16_11_45_1_sva_dfm_1, buf_acc_data_16_12_45_1_sva_dfm_1, buf_acc_data_16_13_45_1_sva_dfm_1,
      buf_acc_data_16_14_45_1_sva_dfm_1, buf_acc_data_16_15_45_1_sva_dfm_1, buf_acc_data_16_16_45_1_sva_dfm_1,
      buf_acc_data_16_17_45_1_sva_dfm_1, buf_acc_data_17_0_45_1_sva_dfm_1, buf_acc_data_17_1_45_1_sva_dfm_1,
      buf_acc_data_17_2_45_1_sva_dfm_1, buf_acc_data_17_3_45_1_sva_dfm_1, buf_acc_data_17_4_45_1_sva_dfm_1,
      buf_acc_data_17_5_45_1_sva_dfm_1, buf_acc_data_17_6_45_1_sva_dfm_1, buf_acc_data_17_7_45_1_sva_dfm_1,
      buf_acc_data_17_8_45_1_sva_dfm_1, buf_acc_data_17_9_45_1_sva_dfm_1, buf_acc_data_17_10_45_1_sva_dfm_1,
      buf_acc_data_17_11_45_1_sva_dfm_1, buf_acc_data_17_12_45_1_sva_dfm_1, buf_acc_data_17_13_45_1_sva_dfm_1,
      buf_acc_data_17_14_45_1_sva_dfm_1, buf_acc_data_17_15_45_1_sva_dfm_1, buf_acc_data_17_16_45_1_sva_dfm_1,
      buf_acc_data_17_17_45_1_sva_dfm_1, {CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_2
      , CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_2
      , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0});
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_56_46_1[10])
      & (~((CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_45_1_1[44:30]==15'b111111111111111)
      & (CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_56_46_1[9:0]==10'b1111111111)));
  assign CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_56_46_1[10])
      | (~((CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_45_1_1[44:30]!=15'b000000000000000)
      | (CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_56_46_1[9:0]!=10'b0000000000))));
  assign CONVOLUTION_LOOP_for_for_for_if_mux_973_nl = MUX_s_1_2_2(buf_acc_data_0_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_980_nl = MUX_s_1_2_2(buf_acc_data_0_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign buf_acc_data_0_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_973_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_980_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_974_nl = MUX_s_1_2_2(buf_acc_data_0_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_982_nl = MUX_s_1_2_2(buf_acc_data_0_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign buf_acc_data_0_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_974_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_982_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_975_nl = MUX_s_1_2_2(buf_acc_data_0_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_984_nl = MUX_s_1_2_2(buf_acc_data_0_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign buf_acc_data_0_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_975_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_984_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_976_nl = MUX_s_1_2_2(buf_acc_data_0_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_986_nl = MUX_s_1_2_2(buf_acc_data_0_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign buf_acc_data_0_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_976_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_986_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_977_nl = MUX_s_1_2_2(buf_acc_data_0_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_988_nl = MUX_s_1_2_2(buf_acc_data_0_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign buf_acc_data_0_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_977_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_988_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_978_nl = MUX_s_1_2_2(buf_acc_data_0_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_990_nl = MUX_s_1_2_2(buf_acc_data_0_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign buf_acc_data_0_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_978_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_990_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_979_nl = MUX_s_1_2_2(buf_acc_data_0_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_992_nl = MUX_s_1_2_2(buf_acc_data_0_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign buf_acc_data_0_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_979_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_992_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_980_nl = MUX_s_1_2_2(buf_acc_data_0_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_994_nl = MUX_s_1_2_2(buf_acc_data_0_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign buf_acc_data_0_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_980_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_994_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_981_nl = MUX_s_1_2_2(buf_acc_data_0_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_996_nl = MUX_s_1_2_2(buf_acc_data_0_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign buf_acc_data_0_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_981_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_996_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_982_nl = MUX_s_1_2_2(buf_acc_data_0_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_998_nl = MUX_s_1_2_2(buf_acc_data_0_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign buf_acc_data_0_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_982_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_998_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_983_nl = MUX_s_1_2_2(buf_acc_data_0_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl = MUX_s_1_2_2(buf_acc_data_0_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign buf_acc_data_0_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_983_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_984_nl = MUX_s_1_2_2(buf_acc_data_0_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl = MUX_s_1_2_2(buf_acc_data_0_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign buf_acc_data_0_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_984_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_985_nl = MUX_s_1_2_2(buf_acc_data_0_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl = MUX_s_1_2_2(buf_acc_data_0_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign buf_acc_data_0_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_985_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_986_nl = MUX_s_1_2_2(buf_acc_data_0_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl = MUX_s_1_2_2(buf_acc_data_0_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign buf_acc_data_0_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_986_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_987_nl = MUX_s_1_2_2(buf_acc_data_0_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl = MUX_s_1_2_2(buf_acc_data_0_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign buf_acc_data_0_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_987_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_988_nl = MUX_s_1_2_2(buf_acc_data_0_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl = MUX_s_1_2_2(buf_acc_data_0_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign buf_acc_data_0_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_988_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_989_nl = MUX_s_1_2_2(buf_acc_data_0_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl = MUX_s_1_2_2(buf_acc_data_0_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign buf_acc_data_0_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_989_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_990_nl = MUX_s_1_2_2(buf_acc_data_0_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl = MUX_s_1_2_2(buf_acc_data_0_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign buf_acc_data_0_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_990_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_991_nl = MUX_s_1_2_2(buf_acc_data_1_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl = MUX_s_1_2_2(buf_acc_data_1_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign buf_acc_data_1_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_991_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_992_nl = MUX_s_1_2_2(buf_acc_data_1_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl = MUX_s_1_2_2(buf_acc_data_1_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign buf_acc_data_1_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_992_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_993_nl = MUX_s_1_2_2(buf_acc_data_1_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl = MUX_s_1_2_2(buf_acc_data_1_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign buf_acc_data_1_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_993_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_994_nl = MUX_s_1_2_2(buf_acc_data_1_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl = MUX_s_1_2_2(buf_acc_data_1_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign buf_acc_data_1_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_994_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_995_nl = MUX_s_1_2_2(buf_acc_data_1_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl = MUX_s_1_2_2(buf_acc_data_1_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign buf_acc_data_1_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_995_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_996_nl = MUX_s_1_2_2(buf_acc_data_1_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl = MUX_s_1_2_2(buf_acc_data_1_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign buf_acc_data_1_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_996_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_997_nl = MUX_s_1_2_2(buf_acc_data_1_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl = MUX_s_1_2_2(buf_acc_data_1_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign buf_acc_data_1_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_997_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_998_nl = MUX_s_1_2_2(buf_acc_data_1_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl = MUX_s_1_2_2(buf_acc_data_1_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign buf_acc_data_1_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_998_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_999_nl = MUX_s_1_2_2(buf_acc_data_1_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl = MUX_s_1_2_2(buf_acc_data_1_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign buf_acc_data_1_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_999_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl = MUX_s_1_2_2(buf_acc_data_1_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl = MUX_s_1_2_2(buf_acc_data_1_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign buf_acc_data_1_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl = MUX_s_1_2_2(buf_acc_data_1_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl = MUX_s_1_2_2(buf_acc_data_1_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign buf_acc_data_1_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl = MUX_s_1_2_2(buf_acc_data_1_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl = MUX_s_1_2_2(buf_acc_data_1_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign buf_acc_data_1_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl = MUX_s_1_2_2(buf_acc_data_1_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl = MUX_s_1_2_2(buf_acc_data_1_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign buf_acc_data_1_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl = MUX_s_1_2_2(buf_acc_data_1_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl = MUX_s_1_2_2(buf_acc_data_1_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign buf_acc_data_1_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl = MUX_s_1_2_2(buf_acc_data_1_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl = MUX_s_1_2_2(buf_acc_data_1_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign buf_acc_data_1_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl = MUX_s_1_2_2(buf_acc_data_1_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl = MUX_s_1_2_2(buf_acc_data_1_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign buf_acc_data_1_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl = MUX_s_1_2_2(buf_acc_data_1_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl = MUX_s_1_2_2(buf_acc_data_1_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign buf_acc_data_1_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl = MUX_s_1_2_2(buf_acc_data_1_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl = MUX_s_1_2_2(buf_acc_data_1_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign buf_acc_data_1_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl = MUX_s_1_2_2(buf_acc_data_2_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl = MUX_s_1_2_2(buf_acc_data_2_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign buf_acc_data_2_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl = MUX_s_1_2_2(buf_acc_data_2_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl = MUX_s_1_2_2(buf_acc_data_2_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign buf_acc_data_2_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl = MUX_s_1_2_2(buf_acc_data_2_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl = MUX_s_1_2_2(buf_acc_data_2_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign buf_acc_data_2_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl = MUX_s_1_2_2(buf_acc_data_2_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl = MUX_s_1_2_2(buf_acc_data_2_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign buf_acc_data_2_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl = MUX_s_1_2_2(buf_acc_data_2_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl = MUX_s_1_2_2(buf_acc_data_2_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign buf_acc_data_2_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl = MUX_s_1_2_2(buf_acc_data_2_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl = MUX_s_1_2_2(buf_acc_data_2_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign buf_acc_data_2_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl = MUX_s_1_2_2(buf_acc_data_2_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl = MUX_s_1_2_2(buf_acc_data_2_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign buf_acc_data_2_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl = MUX_s_1_2_2(buf_acc_data_2_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl = MUX_s_1_2_2(buf_acc_data_2_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign buf_acc_data_2_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl = MUX_s_1_2_2(buf_acc_data_2_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl = MUX_s_1_2_2(buf_acc_data_2_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign buf_acc_data_2_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl = MUX_s_1_2_2(buf_acc_data_2_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl = MUX_s_1_2_2(buf_acc_data_2_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign buf_acc_data_2_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl = MUX_s_1_2_2(buf_acc_data_2_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl = MUX_s_1_2_2(buf_acc_data_2_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign buf_acc_data_2_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl = MUX_s_1_2_2(buf_acc_data_2_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl = MUX_s_1_2_2(buf_acc_data_2_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign buf_acc_data_2_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl = MUX_s_1_2_2(buf_acc_data_2_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl = MUX_s_1_2_2(buf_acc_data_2_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign buf_acc_data_2_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl = MUX_s_1_2_2(buf_acc_data_2_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl = MUX_s_1_2_2(buf_acc_data_2_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign buf_acc_data_2_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl = MUX_s_1_2_2(buf_acc_data_2_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl = MUX_s_1_2_2(buf_acc_data_2_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign buf_acc_data_2_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl = MUX_s_1_2_2(buf_acc_data_2_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl = MUX_s_1_2_2(buf_acc_data_2_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign buf_acc_data_2_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl = MUX_s_1_2_2(buf_acc_data_2_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl = MUX_s_1_2_2(buf_acc_data_2_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign buf_acc_data_2_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl = MUX_s_1_2_2(buf_acc_data_2_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl = MUX_s_1_2_2(buf_acc_data_2_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign buf_acc_data_2_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl = MUX_s_1_2_2(buf_acc_data_3_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl = MUX_s_1_2_2(buf_acc_data_3_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign buf_acc_data_3_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl = MUX_s_1_2_2(buf_acc_data_3_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl = MUX_s_1_2_2(buf_acc_data_3_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign buf_acc_data_3_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl = MUX_s_1_2_2(buf_acc_data_3_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl = MUX_s_1_2_2(buf_acc_data_3_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign buf_acc_data_3_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl = MUX_s_1_2_2(buf_acc_data_3_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl = MUX_s_1_2_2(buf_acc_data_3_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign buf_acc_data_3_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl = MUX_s_1_2_2(buf_acc_data_3_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl = MUX_s_1_2_2(buf_acc_data_3_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign buf_acc_data_3_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl = MUX_s_1_2_2(buf_acc_data_3_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl = MUX_s_1_2_2(buf_acc_data_3_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign buf_acc_data_3_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl = MUX_s_1_2_2(buf_acc_data_3_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl = MUX_s_1_2_2(buf_acc_data_3_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign buf_acc_data_3_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl = MUX_s_1_2_2(buf_acc_data_3_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl = MUX_s_1_2_2(buf_acc_data_3_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign buf_acc_data_3_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl = MUX_s_1_2_2(buf_acc_data_3_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl = MUX_s_1_2_2(buf_acc_data_3_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign buf_acc_data_3_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl = MUX_s_1_2_2(buf_acc_data_3_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl = MUX_s_1_2_2(buf_acc_data_3_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign buf_acc_data_3_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl = MUX_s_1_2_2(buf_acc_data_3_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl = MUX_s_1_2_2(buf_acc_data_3_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign buf_acc_data_3_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl = MUX_s_1_2_2(buf_acc_data_3_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl = MUX_s_1_2_2(buf_acc_data_3_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign buf_acc_data_3_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl = MUX_s_1_2_2(buf_acc_data_3_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl = MUX_s_1_2_2(buf_acc_data_3_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign buf_acc_data_3_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl = MUX_s_1_2_2(buf_acc_data_3_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl = MUX_s_1_2_2(buf_acc_data_3_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign buf_acc_data_3_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl = MUX_s_1_2_2(buf_acc_data_3_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl = MUX_s_1_2_2(buf_acc_data_3_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign buf_acc_data_3_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl = MUX_s_1_2_2(buf_acc_data_3_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl = MUX_s_1_2_2(buf_acc_data_3_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign buf_acc_data_3_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl = MUX_s_1_2_2(buf_acc_data_3_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl = MUX_s_1_2_2(buf_acc_data_3_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign buf_acc_data_3_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl = MUX_s_1_2_2(buf_acc_data_3_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl = MUX_s_1_2_2(buf_acc_data_3_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign buf_acc_data_3_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl = MUX_s_1_2_2(buf_acc_data_4_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl = MUX_s_1_2_2(buf_acc_data_4_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign buf_acc_data_4_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl = MUX_s_1_2_2(buf_acc_data_4_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl = MUX_s_1_2_2(buf_acc_data_4_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign buf_acc_data_4_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl = MUX_s_1_2_2(buf_acc_data_4_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl = MUX_s_1_2_2(buf_acc_data_4_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign buf_acc_data_4_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl = MUX_s_1_2_2(buf_acc_data_4_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl = MUX_s_1_2_2(buf_acc_data_4_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign buf_acc_data_4_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl = MUX_s_1_2_2(buf_acc_data_4_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl = MUX_s_1_2_2(buf_acc_data_4_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign buf_acc_data_4_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl = MUX_s_1_2_2(buf_acc_data_4_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl = MUX_s_1_2_2(buf_acc_data_4_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign buf_acc_data_4_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl = MUX_s_1_2_2(buf_acc_data_4_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl = MUX_s_1_2_2(buf_acc_data_4_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign buf_acc_data_4_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl = MUX_s_1_2_2(buf_acc_data_4_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl = MUX_s_1_2_2(buf_acc_data_4_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign buf_acc_data_4_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl = MUX_s_1_2_2(buf_acc_data_4_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl = MUX_s_1_2_2(buf_acc_data_4_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign buf_acc_data_4_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl = MUX_s_1_2_2(buf_acc_data_4_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl = MUX_s_1_2_2(buf_acc_data_4_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign buf_acc_data_4_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl = MUX_s_1_2_2(buf_acc_data_4_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl = MUX_s_1_2_2(buf_acc_data_4_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign buf_acc_data_4_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl = MUX_s_1_2_2(buf_acc_data_4_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl = MUX_s_1_2_2(buf_acc_data_4_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign buf_acc_data_4_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl = MUX_s_1_2_2(buf_acc_data_4_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl = MUX_s_1_2_2(buf_acc_data_4_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign buf_acc_data_4_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl = MUX_s_1_2_2(buf_acc_data_4_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl = MUX_s_1_2_2(buf_acc_data_4_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign buf_acc_data_4_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl = MUX_s_1_2_2(buf_acc_data_4_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl = MUX_s_1_2_2(buf_acc_data_4_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign buf_acc_data_4_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl = MUX_s_1_2_2(buf_acc_data_4_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl = MUX_s_1_2_2(buf_acc_data_4_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign buf_acc_data_4_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl = MUX_s_1_2_2(buf_acc_data_4_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl = MUX_s_1_2_2(buf_acc_data_4_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign buf_acc_data_4_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl = MUX_s_1_2_2(buf_acc_data_4_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl = MUX_s_1_2_2(buf_acc_data_4_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign buf_acc_data_4_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl = MUX_s_1_2_2(buf_acc_data_5_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl = MUX_s_1_2_2(buf_acc_data_5_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign buf_acc_data_5_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl = MUX_s_1_2_2(buf_acc_data_5_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl = MUX_s_1_2_2(buf_acc_data_5_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign buf_acc_data_5_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl = MUX_s_1_2_2(buf_acc_data_5_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl = MUX_s_1_2_2(buf_acc_data_5_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign buf_acc_data_5_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl = MUX_s_1_2_2(buf_acc_data_5_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl = MUX_s_1_2_2(buf_acc_data_5_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign buf_acc_data_5_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl = MUX_s_1_2_2(buf_acc_data_5_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl = MUX_s_1_2_2(buf_acc_data_5_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign buf_acc_data_5_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl = MUX_s_1_2_2(buf_acc_data_5_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl = MUX_s_1_2_2(buf_acc_data_5_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign buf_acc_data_5_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl = MUX_s_1_2_2(buf_acc_data_5_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl = MUX_s_1_2_2(buf_acc_data_5_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign buf_acc_data_5_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl = MUX_s_1_2_2(buf_acc_data_5_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl = MUX_s_1_2_2(buf_acc_data_5_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign buf_acc_data_5_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl = MUX_s_1_2_2(buf_acc_data_5_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl = MUX_s_1_2_2(buf_acc_data_5_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign buf_acc_data_5_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl = MUX_s_1_2_2(buf_acc_data_5_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl = MUX_s_1_2_2(buf_acc_data_5_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign buf_acc_data_5_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl = MUX_s_1_2_2(buf_acc_data_5_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl = MUX_s_1_2_2(buf_acc_data_5_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign buf_acc_data_5_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl = MUX_s_1_2_2(buf_acc_data_5_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl = MUX_s_1_2_2(buf_acc_data_5_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign buf_acc_data_5_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl = MUX_s_1_2_2(buf_acc_data_5_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl = MUX_s_1_2_2(buf_acc_data_5_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign buf_acc_data_5_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl = MUX_s_1_2_2(buf_acc_data_5_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl = MUX_s_1_2_2(buf_acc_data_5_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign buf_acc_data_5_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl = MUX_s_1_2_2(buf_acc_data_5_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl = MUX_s_1_2_2(buf_acc_data_5_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign buf_acc_data_5_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl = MUX_s_1_2_2(buf_acc_data_5_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl = MUX_s_1_2_2(buf_acc_data_5_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign buf_acc_data_5_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl = MUX_s_1_2_2(buf_acc_data_5_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl = MUX_s_1_2_2(buf_acc_data_5_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign buf_acc_data_5_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl = MUX_s_1_2_2(buf_acc_data_5_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl = MUX_s_1_2_2(buf_acc_data_5_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign buf_acc_data_5_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl = MUX_s_1_2_2(buf_acc_data_6_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl = MUX_s_1_2_2(buf_acc_data_6_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign buf_acc_data_6_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl = MUX_s_1_2_2(buf_acc_data_6_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl = MUX_s_1_2_2(buf_acc_data_6_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign buf_acc_data_6_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl = MUX_s_1_2_2(buf_acc_data_6_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl = MUX_s_1_2_2(buf_acc_data_6_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign buf_acc_data_6_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl = MUX_s_1_2_2(buf_acc_data_6_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl = MUX_s_1_2_2(buf_acc_data_6_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign buf_acc_data_6_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl = MUX_s_1_2_2(buf_acc_data_6_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl = MUX_s_1_2_2(buf_acc_data_6_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign buf_acc_data_6_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl = MUX_s_1_2_2(buf_acc_data_6_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl = MUX_s_1_2_2(buf_acc_data_6_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign buf_acc_data_6_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl = MUX_s_1_2_2(buf_acc_data_6_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl = MUX_s_1_2_2(buf_acc_data_6_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign buf_acc_data_6_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl = MUX_s_1_2_2(buf_acc_data_6_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl = MUX_s_1_2_2(buf_acc_data_6_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign buf_acc_data_6_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl = MUX_s_1_2_2(buf_acc_data_6_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl = MUX_s_1_2_2(buf_acc_data_6_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign buf_acc_data_6_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl = MUX_s_1_2_2(buf_acc_data_6_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl = MUX_s_1_2_2(buf_acc_data_6_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign buf_acc_data_6_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl = MUX_s_1_2_2(buf_acc_data_6_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl = MUX_s_1_2_2(buf_acc_data_6_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign buf_acc_data_6_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl = MUX_s_1_2_2(buf_acc_data_6_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl = MUX_s_1_2_2(buf_acc_data_6_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign buf_acc_data_6_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl = MUX_s_1_2_2(buf_acc_data_6_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl = MUX_s_1_2_2(buf_acc_data_6_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign buf_acc_data_6_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl = MUX_s_1_2_2(buf_acc_data_6_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl = MUX_s_1_2_2(buf_acc_data_6_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign buf_acc_data_6_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl = MUX_s_1_2_2(buf_acc_data_6_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl = MUX_s_1_2_2(buf_acc_data_6_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign buf_acc_data_6_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl = MUX_s_1_2_2(buf_acc_data_6_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl = MUX_s_1_2_2(buf_acc_data_6_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign buf_acc_data_6_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl = MUX_s_1_2_2(buf_acc_data_6_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl = MUX_s_1_2_2(buf_acc_data_6_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign buf_acc_data_6_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl = MUX_s_1_2_2(buf_acc_data_6_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl = MUX_s_1_2_2(buf_acc_data_6_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign buf_acc_data_6_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl = MUX_s_1_2_2(buf_acc_data_7_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl = MUX_s_1_2_2(buf_acc_data_7_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign buf_acc_data_7_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl = MUX_s_1_2_2(buf_acc_data_7_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl = MUX_s_1_2_2(buf_acc_data_7_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign buf_acc_data_7_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl = MUX_s_1_2_2(buf_acc_data_7_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl = MUX_s_1_2_2(buf_acc_data_7_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign buf_acc_data_7_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl = MUX_s_1_2_2(buf_acc_data_7_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl = MUX_s_1_2_2(buf_acc_data_7_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign buf_acc_data_7_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl = MUX_s_1_2_2(buf_acc_data_7_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl = MUX_s_1_2_2(buf_acc_data_7_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign buf_acc_data_7_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl = MUX_s_1_2_2(buf_acc_data_7_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl = MUX_s_1_2_2(buf_acc_data_7_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign buf_acc_data_7_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl = MUX_s_1_2_2(buf_acc_data_7_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl = MUX_s_1_2_2(buf_acc_data_7_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign buf_acc_data_7_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl = MUX_s_1_2_2(buf_acc_data_7_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl = MUX_s_1_2_2(buf_acc_data_7_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign buf_acc_data_7_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl = MUX_s_1_2_2(buf_acc_data_7_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl = MUX_s_1_2_2(buf_acc_data_7_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign buf_acc_data_7_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl = MUX_s_1_2_2(buf_acc_data_7_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl = MUX_s_1_2_2(buf_acc_data_7_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign buf_acc_data_7_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl = MUX_s_1_2_2(buf_acc_data_7_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl = MUX_s_1_2_2(buf_acc_data_7_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign buf_acc_data_7_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl = MUX_s_1_2_2(buf_acc_data_7_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl = MUX_s_1_2_2(buf_acc_data_7_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign buf_acc_data_7_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl = MUX_s_1_2_2(buf_acc_data_7_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl = MUX_s_1_2_2(buf_acc_data_7_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1);
  assign buf_acc_data_7_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl = MUX_s_1_2_2(buf_acc_data_7_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl = MUX_s_1_2_2(buf_acc_data_7_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1);
  assign buf_acc_data_7_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl = MUX_s_1_2_2(buf_acc_data_7_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl = MUX_s_1_2_2(buf_acc_data_7_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1);
  assign buf_acc_data_7_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl = MUX_s_1_2_2(buf_acc_data_7_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl = MUX_s_1_2_2(buf_acc_data_7_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1);
  assign buf_acc_data_7_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl = MUX_s_1_2_2(buf_acc_data_7_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl = MUX_s_1_2_2(buf_acc_data_7_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1);
  assign buf_acc_data_7_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl = MUX_s_1_2_2(buf_acc_data_7_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl = MUX_s_1_2_2(buf_acc_data_7_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1);
  assign buf_acc_data_7_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl = MUX_s_1_2_2(buf_acc_data_8_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl = MUX_s_1_2_2(buf_acc_data_8_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1);
  assign buf_acc_data_8_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl = MUX_s_1_2_2(buf_acc_data_8_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl = MUX_s_1_2_2(buf_acc_data_8_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1);
  assign buf_acc_data_8_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl = MUX_s_1_2_2(buf_acc_data_8_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl = MUX_s_1_2_2(buf_acc_data_8_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1);
  assign buf_acc_data_8_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl = MUX_s_1_2_2(buf_acc_data_8_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl = MUX_s_1_2_2(buf_acc_data_8_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1);
  assign buf_acc_data_8_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl = MUX_s_1_2_2(buf_acc_data_8_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl = MUX_s_1_2_2(buf_acc_data_8_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1);
  assign buf_acc_data_8_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl = MUX_s_1_2_2(buf_acc_data_8_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl = MUX_s_1_2_2(buf_acc_data_8_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1);
  assign buf_acc_data_8_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl = MUX_s_1_2_2(buf_acc_data_8_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl = MUX_s_1_2_2(buf_acc_data_8_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1);
  assign buf_acc_data_8_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl = MUX_s_1_2_2(buf_acc_data_8_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl = MUX_s_1_2_2(buf_acc_data_8_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1);
  assign buf_acc_data_8_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl = MUX_s_1_2_2(buf_acc_data_8_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl = MUX_s_1_2_2(buf_acc_data_8_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1);
  assign buf_acc_data_8_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl = MUX_s_1_2_2(buf_acc_data_8_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl = MUX_s_1_2_2(buf_acc_data_8_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1);
  assign buf_acc_data_8_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl = MUX_s_1_2_2(buf_acc_data_8_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl = MUX_s_1_2_2(buf_acc_data_8_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1);
  assign buf_acc_data_8_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl = MUX_s_1_2_2(buf_acc_data_8_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl = MUX_s_1_2_2(buf_acc_data_8_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1);
  assign buf_acc_data_8_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl = MUX_s_1_2_2(buf_acc_data_8_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl = MUX_s_1_2_2(buf_acc_data_8_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1);
  assign buf_acc_data_8_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl = MUX_s_1_2_2(buf_acc_data_8_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl = MUX_s_1_2_2(buf_acc_data_8_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1);
  assign buf_acc_data_8_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl = MUX_s_1_2_2(buf_acc_data_8_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl = MUX_s_1_2_2(buf_acc_data_8_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1);
  assign buf_acc_data_8_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl = MUX_s_1_2_2(buf_acc_data_8_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl = MUX_s_1_2_2(buf_acc_data_8_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1);
  assign buf_acc_data_8_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl = MUX_s_1_2_2(buf_acc_data_8_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl = MUX_s_1_2_2(buf_acc_data_8_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1);
  assign buf_acc_data_8_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl = MUX_s_1_2_2(buf_acc_data_8_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl = MUX_s_1_2_2(buf_acc_data_8_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1);
  assign buf_acc_data_8_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl = MUX_s_1_2_2(buf_acc_data_9_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl = MUX_s_1_2_2(buf_acc_data_9_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1);
  assign buf_acc_data_9_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl = MUX_s_1_2_2(buf_acc_data_9_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl = MUX_s_1_2_2(buf_acc_data_9_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1);
  assign buf_acc_data_9_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl = MUX_s_1_2_2(buf_acc_data_9_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl = MUX_s_1_2_2(buf_acc_data_9_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1);
  assign buf_acc_data_9_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl = MUX_s_1_2_2(buf_acc_data_9_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl = MUX_s_1_2_2(buf_acc_data_9_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1);
  assign buf_acc_data_9_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl = MUX_s_1_2_2(buf_acc_data_9_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl = MUX_s_1_2_2(buf_acc_data_9_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1);
  assign buf_acc_data_9_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl = MUX_s_1_2_2(buf_acc_data_9_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl = MUX_s_1_2_2(buf_acc_data_9_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1);
  assign buf_acc_data_9_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl = MUX_s_1_2_2(buf_acc_data_9_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl = MUX_s_1_2_2(buf_acc_data_9_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1);
  assign buf_acc_data_9_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl = MUX_s_1_2_2(buf_acc_data_9_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl = MUX_s_1_2_2(buf_acc_data_9_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1);
  assign buf_acc_data_9_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl = MUX_s_1_2_2(buf_acc_data_9_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl = MUX_s_1_2_2(buf_acc_data_9_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1);
  assign buf_acc_data_9_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl = MUX_s_1_2_2(buf_acc_data_9_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl = MUX_s_1_2_2(buf_acc_data_9_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1);
  assign buf_acc_data_9_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl = MUX_s_1_2_2(buf_acc_data_9_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl = MUX_s_1_2_2(buf_acc_data_9_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1);
  assign buf_acc_data_9_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl = MUX_s_1_2_2(buf_acc_data_9_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl = MUX_s_1_2_2(buf_acc_data_9_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1);
  assign buf_acc_data_9_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl = MUX_s_1_2_2(buf_acc_data_9_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl = MUX_s_1_2_2(buf_acc_data_9_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1);
  assign buf_acc_data_9_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl = MUX_s_1_2_2(buf_acc_data_9_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl = MUX_s_1_2_2(buf_acc_data_9_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1);
  assign buf_acc_data_9_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl = MUX_s_1_2_2(buf_acc_data_9_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl = MUX_s_1_2_2(buf_acc_data_9_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1);
  assign buf_acc_data_9_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl = MUX_s_1_2_2(buf_acc_data_9_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl = MUX_s_1_2_2(buf_acc_data_9_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1);
  assign buf_acc_data_9_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl = MUX_s_1_2_2(buf_acc_data_9_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl = MUX_s_1_2_2(buf_acc_data_9_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1);
  assign buf_acc_data_9_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl = MUX_s_1_2_2(buf_acc_data_9_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl = MUX_s_1_2_2(buf_acc_data_9_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1);
  assign buf_acc_data_9_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl = MUX_s_1_2_2(buf_acc_data_10_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl = MUX_s_1_2_2(buf_acc_data_10_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1);
  assign buf_acc_data_10_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl = MUX_s_1_2_2(buf_acc_data_10_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl = MUX_s_1_2_2(buf_acc_data_10_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1);
  assign buf_acc_data_10_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl = MUX_s_1_2_2(buf_acc_data_10_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl = MUX_s_1_2_2(buf_acc_data_10_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1);
  assign buf_acc_data_10_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl = MUX_s_1_2_2(buf_acc_data_10_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl = MUX_s_1_2_2(buf_acc_data_10_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1);
  assign buf_acc_data_10_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl = MUX_s_1_2_2(buf_acc_data_10_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl = MUX_s_1_2_2(buf_acc_data_10_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1);
  assign buf_acc_data_10_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl = MUX_s_1_2_2(buf_acc_data_10_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl = MUX_s_1_2_2(buf_acc_data_10_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1);
  assign buf_acc_data_10_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl = MUX_s_1_2_2(buf_acc_data_10_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl = MUX_s_1_2_2(buf_acc_data_10_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign buf_acc_data_10_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl = MUX_s_1_2_2(buf_acc_data_10_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl = MUX_s_1_2_2(buf_acc_data_10_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign buf_acc_data_10_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl = MUX_s_1_2_2(buf_acc_data_10_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl = MUX_s_1_2_2(buf_acc_data_10_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign buf_acc_data_10_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl = MUX_s_1_2_2(buf_acc_data_10_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl = MUX_s_1_2_2(buf_acc_data_10_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign buf_acc_data_10_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl = MUX_s_1_2_2(buf_acc_data_10_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl = MUX_s_1_2_2(buf_acc_data_10_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign buf_acc_data_10_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl = MUX_s_1_2_2(buf_acc_data_10_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl = MUX_s_1_2_2(buf_acc_data_10_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign buf_acc_data_10_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl = MUX_s_1_2_2(buf_acc_data_10_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl = MUX_s_1_2_2(buf_acc_data_10_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign buf_acc_data_10_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl = MUX_s_1_2_2(buf_acc_data_10_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl = MUX_s_1_2_2(buf_acc_data_10_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign buf_acc_data_10_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl = MUX_s_1_2_2(buf_acc_data_10_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl = MUX_s_1_2_2(buf_acc_data_10_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign buf_acc_data_10_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl = MUX_s_1_2_2(buf_acc_data_10_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl = MUX_s_1_2_2(buf_acc_data_10_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign buf_acc_data_10_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl = MUX_s_1_2_2(buf_acc_data_10_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl = MUX_s_1_2_2(buf_acc_data_10_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign buf_acc_data_10_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl = MUX_s_1_2_2(buf_acc_data_10_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl = MUX_s_1_2_2(buf_acc_data_10_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign buf_acc_data_10_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl = MUX_s_1_2_2(buf_acc_data_11_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl = MUX_s_1_2_2(buf_acc_data_11_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign buf_acc_data_11_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl = MUX_s_1_2_2(buf_acc_data_11_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl = MUX_s_1_2_2(buf_acc_data_11_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign buf_acc_data_11_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl = MUX_s_1_2_2(buf_acc_data_11_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl = MUX_s_1_2_2(buf_acc_data_11_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign buf_acc_data_11_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl = MUX_s_1_2_2(buf_acc_data_11_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl = MUX_s_1_2_2(buf_acc_data_11_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign buf_acc_data_11_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl = MUX_s_1_2_2(buf_acc_data_11_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl = MUX_s_1_2_2(buf_acc_data_11_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign buf_acc_data_11_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl = MUX_s_1_2_2(buf_acc_data_11_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl = MUX_s_1_2_2(buf_acc_data_11_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign buf_acc_data_11_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl = MUX_s_1_2_2(buf_acc_data_11_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl = MUX_s_1_2_2(buf_acc_data_11_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign buf_acc_data_11_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl = MUX_s_1_2_2(buf_acc_data_11_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl = MUX_s_1_2_2(buf_acc_data_11_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign buf_acc_data_11_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl = MUX_s_1_2_2(buf_acc_data_11_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl = MUX_s_1_2_2(buf_acc_data_11_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign buf_acc_data_11_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl = MUX_s_1_2_2(buf_acc_data_11_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl = MUX_s_1_2_2(buf_acc_data_11_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign buf_acc_data_11_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl = MUX_s_1_2_2(buf_acc_data_11_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl = MUX_s_1_2_2(buf_acc_data_11_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign buf_acc_data_11_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl = MUX_s_1_2_2(buf_acc_data_11_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl = MUX_s_1_2_2(buf_acc_data_11_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign buf_acc_data_11_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl = MUX_s_1_2_2(buf_acc_data_11_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl = MUX_s_1_2_2(buf_acc_data_11_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign buf_acc_data_11_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl = MUX_s_1_2_2(buf_acc_data_11_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl = MUX_s_1_2_2(buf_acc_data_11_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign buf_acc_data_11_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl = MUX_s_1_2_2(buf_acc_data_11_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl = MUX_s_1_2_2(buf_acc_data_11_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign buf_acc_data_11_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl = MUX_s_1_2_2(buf_acc_data_11_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl = MUX_s_1_2_2(buf_acc_data_11_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign buf_acc_data_11_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl = MUX_s_1_2_2(buf_acc_data_11_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl = MUX_s_1_2_2(buf_acc_data_11_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign buf_acc_data_11_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl = MUX_s_1_2_2(buf_acc_data_11_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl = MUX_s_1_2_2(buf_acc_data_11_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign buf_acc_data_11_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl = MUX_s_1_2_2(buf_acc_data_12_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl = MUX_s_1_2_2(buf_acc_data_12_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign buf_acc_data_12_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl = MUX_s_1_2_2(buf_acc_data_12_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl = MUX_s_1_2_2(buf_acc_data_12_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign buf_acc_data_12_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl = MUX_s_1_2_2(buf_acc_data_12_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl = MUX_s_1_2_2(buf_acc_data_12_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign buf_acc_data_12_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl = MUX_s_1_2_2(buf_acc_data_12_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl = MUX_s_1_2_2(buf_acc_data_12_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign buf_acc_data_12_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl = MUX_s_1_2_2(buf_acc_data_12_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl = MUX_s_1_2_2(buf_acc_data_12_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign buf_acc_data_12_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl = MUX_s_1_2_2(buf_acc_data_12_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl = MUX_s_1_2_2(buf_acc_data_12_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign buf_acc_data_12_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl = MUX_s_1_2_2(buf_acc_data_12_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl = MUX_s_1_2_2(buf_acc_data_12_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign buf_acc_data_12_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl = MUX_s_1_2_2(buf_acc_data_12_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl = MUX_s_1_2_2(buf_acc_data_12_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign buf_acc_data_12_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl = MUX_s_1_2_2(buf_acc_data_12_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl = MUX_s_1_2_2(buf_acc_data_12_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign buf_acc_data_12_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl = MUX_s_1_2_2(buf_acc_data_12_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl = MUX_s_1_2_2(buf_acc_data_12_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign buf_acc_data_12_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl = MUX_s_1_2_2(buf_acc_data_12_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl = MUX_s_1_2_2(buf_acc_data_12_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign buf_acc_data_12_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl = MUX_s_1_2_2(buf_acc_data_12_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl = MUX_s_1_2_2(buf_acc_data_12_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign buf_acc_data_12_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl = MUX_s_1_2_2(buf_acc_data_12_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl = MUX_s_1_2_2(buf_acc_data_12_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign buf_acc_data_12_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl = MUX_s_1_2_2(buf_acc_data_12_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl = MUX_s_1_2_2(buf_acc_data_12_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign buf_acc_data_12_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl = MUX_s_1_2_2(buf_acc_data_12_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl = MUX_s_1_2_2(buf_acc_data_12_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign buf_acc_data_12_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl = MUX_s_1_2_2(buf_acc_data_12_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl = MUX_s_1_2_2(buf_acc_data_12_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign buf_acc_data_12_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl = MUX_s_1_2_2(buf_acc_data_12_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl = MUX_s_1_2_2(buf_acc_data_12_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign buf_acc_data_12_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl = MUX_s_1_2_2(buf_acc_data_12_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl = MUX_s_1_2_2(buf_acc_data_12_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign buf_acc_data_12_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl = MUX_s_1_2_2(buf_acc_data_13_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl = MUX_s_1_2_2(buf_acc_data_13_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign buf_acc_data_13_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl = MUX_s_1_2_2(buf_acc_data_13_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl = MUX_s_1_2_2(buf_acc_data_13_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign buf_acc_data_13_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl = MUX_s_1_2_2(buf_acc_data_13_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl = MUX_s_1_2_2(buf_acc_data_13_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign buf_acc_data_13_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl = MUX_s_1_2_2(buf_acc_data_13_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl = MUX_s_1_2_2(buf_acc_data_13_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign buf_acc_data_13_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl = MUX_s_1_2_2(buf_acc_data_13_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl = MUX_s_1_2_2(buf_acc_data_13_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign buf_acc_data_13_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl = MUX_s_1_2_2(buf_acc_data_13_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl = MUX_s_1_2_2(buf_acc_data_13_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign buf_acc_data_13_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl = MUX_s_1_2_2(buf_acc_data_13_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl = MUX_s_1_2_2(buf_acc_data_13_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign buf_acc_data_13_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl = MUX_s_1_2_2(buf_acc_data_13_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl = MUX_s_1_2_2(buf_acc_data_13_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign buf_acc_data_13_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl = MUX_s_1_2_2(buf_acc_data_13_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl = MUX_s_1_2_2(buf_acc_data_13_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign buf_acc_data_13_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl = MUX_s_1_2_2(buf_acc_data_13_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl = MUX_s_1_2_2(buf_acc_data_13_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign buf_acc_data_13_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl = MUX_s_1_2_2(buf_acc_data_13_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl = MUX_s_1_2_2(buf_acc_data_13_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign buf_acc_data_13_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl = MUX_s_1_2_2(buf_acc_data_13_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl = MUX_s_1_2_2(buf_acc_data_13_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign buf_acc_data_13_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl = MUX_s_1_2_2(buf_acc_data_13_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl = MUX_s_1_2_2(buf_acc_data_13_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign buf_acc_data_13_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl = MUX_s_1_2_2(buf_acc_data_13_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl = MUX_s_1_2_2(buf_acc_data_13_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign buf_acc_data_13_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl = MUX_s_1_2_2(buf_acc_data_13_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl = MUX_s_1_2_2(buf_acc_data_13_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign buf_acc_data_13_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl = MUX_s_1_2_2(buf_acc_data_13_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl = MUX_s_1_2_2(buf_acc_data_13_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign buf_acc_data_13_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl = MUX_s_1_2_2(buf_acc_data_13_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl = MUX_s_1_2_2(buf_acc_data_13_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign buf_acc_data_13_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl = MUX_s_1_2_2(buf_acc_data_13_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl = MUX_s_1_2_2(buf_acc_data_13_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign buf_acc_data_13_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl = MUX_s_1_2_2(buf_acc_data_14_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl = MUX_s_1_2_2(buf_acc_data_14_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign buf_acc_data_14_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl = MUX_s_1_2_2(buf_acc_data_14_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl = MUX_s_1_2_2(buf_acc_data_14_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign buf_acc_data_14_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl = MUX_s_1_2_2(buf_acc_data_14_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl = MUX_s_1_2_2(buf_acc_data_14_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign buf_acc_data_14_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl = MUX_s_1_2_2(buf_acc_data_14_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl = MUX_s_1_2_2(buf_acc_data_14_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign buf_acc_data_14_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl = MUX_s_1_2_2(buf_acc_data_14_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl = MUX_s_1_2_2(buf_acc_data_14_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign buf_acc_data_14_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl = MUX_s_1_2_2(buf_acc_data_14_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl = MUX_s_1_2_2(buf_acc_data_14_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign buf_acc_data_14_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl = MUX_s_1_2_2(buf_acc_data_14_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl = MUX_s_1_2_2(buf_acc_data_14_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign buf_acc_data_14_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl = MUX_s_1_2_2(buf_acc_data_14_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl = MUX_s_1_2_2(buf_acc_data_14_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign buf_acc_data_14_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl = MUX_s_1_2_2(buf_acc_data_14_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl = MUX_s_1_2_2(buf_acc_data_14_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign buf_acc_data_14_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl = MUX_s_1_2_2(buf_acc_data_14_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl = MUX_s_1_2_2(buf_acc_data_14_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign buf_acc_data_14_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl = MUX_s_1_2_2(buf_acc_data_14_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl = MUX_s_1_2_2(buf_acc_data_14_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign buf_acc_data_14_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl = MUX_s_1_2_2(buf_acc_data_14_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl = MUX_s_1_2_2(buf_acc_data_14_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign buf_acc_data_14_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl = MUX_s_1_2_2(buf_acc_data_14_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl = MUX_s_1_2_2(buf_acc_data_14_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign buf_acc_data_14_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl = MUX_s_1_2_2(buf_acc_data_14_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl = MUX_s_1_2_2(buf_acc_data_14_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign buf_acc_data_14_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl = MUX_s_1_2_2(buf_acc_data_14_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl = MUX_s_1_2_2(buf_acc_data_14_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign buf_acc_data_14_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl = MUX_s_1_2_2(buf_acc_data_14_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl = MUX_s_1_2_2(buf_acc_data_14_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign buf_acc_data_14_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl = MUX_s_1_2_2(buf_acc_data_14_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl = MUX_s_1_2_2(buf_acc_data_14_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign buf_acc_data_14_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl = MUX_s_1_2_2(buf_acc_data_14_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl = MUX_s_1_2_2(buf_acc_data_14_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign buf_acc_data_14_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl = MUX_s_1_2_2(buf_acc_data_15_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl = MUX_s_1_2_2(buf_acc_data_15_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign buf_acc_data_15_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl = MUX_s_1_2_2(buf_acc_data_15_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl = MUX_s_1_2_2(buf_acc_data_15_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign buf_acc_data_15_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl = MUX_s_1_2_2(buf_acc_data_15_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl = MUX_s_1_2_2(buf_acc_data_15_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign buf_acc_data_15_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl = MUX_s_1_2_2(buf_acc_data_15_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl = MUX_s_1_2_2(buf_acc_data_15_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign buf_acc_data_15_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl = MUX_s_1_2_2(buf_acc_data_15_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl = MUX_s_1_2_2(buf_acc_data_15_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign buf_acc_data_15_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl = MUX_s_1_2_2(buf_acc_data_15_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl = MUX_s_1_2_2(buf_acc_data_15_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign buf_acc_data_15_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl = MUX_s_1_2_2(buf_acc_data_15_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl = MUX_s_1_2_2(buf_acc_data_15_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign buf_acc_data_15_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl = MUX_s_1_2_2(buf_acc_data_15_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl = MUX_s_1_2_2(buf_acc_data_15_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign buf_acc_data_15_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl = MUX_s_1_2_2(buf_acc_data_15_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl = MUX_s_1_2_2(buf_acc_data_15_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign buf_acc_data_15_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl = MUX_s_1_2_2(buf_acc_data_15_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl = MUX_s_1_2_2(buf_acc_data_15_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign buf_acc_data_15_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl = MUX_s_1_2_2(buf_acc_data_15_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl = MUX_s_1_2_2(buf_acc_data_15_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign buf_acc_data_15_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl = MUX_s_1_2_2(buf_acc_data_15_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl = MUX_s_1_2_2(buf_acc_data_15_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign buf_acc_data_15_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl = MUX_s_1_2_2(buf_acc_data_15_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl = MUX_s_1_2_2(buf_acc_data_15_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign buf_acc_data_15_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl = MUX_s_1_2_2(buf_acc_data_15_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl = MUX_s_1_2_2(buf_acc_data_15_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign buf_acc_data_15_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl = MUX_s_1_2_2(buf_acc_data_15_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl = MUX_s_1_2_2(buf_acc_data_15_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign buf_acc_data_15_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl = MUX_s_1_2_2(buf_acc_data_15_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl = MUX_s_1_2_2(buf_acc_data_15_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign buf_acc_data_15_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl = MUX_s_1_2_2(buf_acc_data_15_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl = MUX_s_1_2_2(buf_acc_data_15_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign buf_acc_data_15_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl = MUX_s_1_2_2(buf_acc_data_15_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl = MUX_s_1_2_2(buf_acc_data_15_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign buf_acc_data_15_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl = MUX_s_1_2_2(buf_acc_data_16_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl = MUX_s_1_2_2(buf_acc_data_16_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign buf_acc_data_16_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl = MUX_s_1_2_2(buf_acc_data_16_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl = MUX_s_1_2_2(buf_acc_data_16_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign buf_acc_data_16_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl = MUX_s_1_2_2(buf_acc_data_16_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl = MUX_s_1_2_2(buf_acc_data_16_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign buf_acc_data_16_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl = MUX_s_1_2_2(buf_acc_data_16_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl = MUX_s_1_2_2(buf_acc_data_16_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign buf_acc_data_16_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl = MUX_s_1_2_2(buf_acc_data_16_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl = MUX_s_1_2_2(buf_acc_data_16_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign buf_acc_data_16_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl = MUX_s_1_2_2(buf_acc_data_16_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl = MUX_s_1_2_2(buf_acc_data_16_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign buf_acc_data_16_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl = MUX_s_1_2_2(buf_acc_data_16_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl = MUX_s_1_2_2(buf_acc_data_16_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign buf_acc_data_16_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl = MUX_s_1_2_2(buf_acc_data_16_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl = MUX_s_1_2_2(buf_acc_data_16_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign buf_acc_data_16_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl = MUX_s_1_2_2(buf_acc_data_16_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl = MUX_s_1_2_2(buf_acc_data_16_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign buf_acc_data_16_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl = MUX_s_1_2_2(buf_acc_data_16_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl = MUX_s_1_2_2(buf_acc_data_16_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign buf_acc_data_16_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl = MUX_s_1_2_2(buf_acc_data_16_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl = MUX_s_1_2_2(buf_acc_data_16_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign buf_acc_data_16_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl = MUX_s_1_2_2(buf_acc_data_16_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl = MUX_s_1_2_2(buf_acc_data_16_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign buf_acc_data_16_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl = MUX_s_1_2_2(buf_acc_data_16_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl = MUX_s_1_2_2(buf_acc_data_16_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign buf_acc_data_16_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl = MUX_s_1_2_2(buf_acc_data_16_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl = MUX_s_1_2_2(buf_acc_data_16_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign buf_acc_data_16_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl = MUX_s_1_2_2(buf_acc_data_16_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl = MUX_s_1_2_2(buf_acc_data_16_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign buf_acc_data_16_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl = MUX_s_1_2_2(buf_acc_data_16_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl = MUX_s_1_2_2(buf_acc_data_16_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign buf_acc_data_16_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl = MUX_s_1_2_2(buf_acc_data_16_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl = MUX_s_1_2_2(buf_acc_data_16_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign buf_acc_data_16_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl = MUX_s_1_2_2(buf_acc_data_16_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl = MUX_s_1_2_2(buf_acc_data_16_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign buf_acc_data_16_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl = MUX_s_1_2_2(buf_acc_data_17_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl = MUX_s_1_2_2(buf_acc_data_17_0_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign buf_acc_data_17_0_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl = MUX_s_1_2_2(buf_acc_data_17_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl = MUX_s_1_2_2(buf_acc_data_17_1_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign buf_acc_data_17_1_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl = MUX_s_1_2_2(buf_acc_data_17_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl = MUX_s_1_2_2(buf_acc_data_17_2_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign buf_acc_data_17_2_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl = MUX_s_1_2_2(buf_acc_data_17_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl = MUX_s_1_2_2(buf_acc_data_17_3_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign buf_acc_data_17_3_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl = MUX_s_1_2_2(buf_acc_data_17_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl = MUX_s_1_2_2(buf_acc_data_17_4_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign buf_acc_data_17_4_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl = MUX_s_1_2_2(buf_acc_data_17_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl = MUX_s_1_2_2(buf_acc_data_17_5_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign buf_acc_data_17_5_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl = MUX_s_1_2_2(buf_acc_data_17_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl = MUX_s_1_2_2(buf_acc_data_17_6_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign buf_acc_data_17_6_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl = MUX_s_1_2_2(buf_acc_data_17_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl = MUX_s_1_2_2(buf_acc_data_17_7_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign buf_acc_data_17_7_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl = MUX_s_1_2_2(buf_acc_data_17_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl = MUX_s_1_2_2(buf_acc_data_17_8_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign buf_acc_data_17_8_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl = MUX_s_1_2_2(buf_acc_data_17_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl = MUX_s_1_2_2(buf_acc_data_17_9_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign buf_acc_data_17_9_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl = MUX_s_1_2_2(buf_acc_data_17_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl = MUX_s_1_2_2(buf_acc_data_17_10_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign buf_acc_data_17_10_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl = MUX_s_1_2_2(buf_acc_data_17_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl = MUX_s_1_2_2(buf_acc_data_17_11_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign buf_acc_data_17_11_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl = MUX_s_1_2_2(buf_acc_data_17_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl = MUX_s_1_2_2(buf_acc_data_17_12_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign buf_acc_data_17_12_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl = MUX_s_1_2_2(buf_acc_data_17_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl = MUX_s_1_2_2(buf_acc_data_17_13_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign buf_acc_data_17_13_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl = MUX_s_1_2_2(buf_acc_data_17_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl = MUX_s_1_2_2(buf_acc_data_17_14_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign buf_acc_data_17_14_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl = MUX_s_1_2_2(buf_acc_data_17_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl = MUX_s_1_2_2(buf_acc_data_17_15_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign buf_acc_data_17_15_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl = MUX_s_1_2_2(buf_acc_data_17_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl = MUX_s_1_2_2(buf_acc_data_17_16_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign buf_acc_data_17_16_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl = MUX_s_1_2_2(buf_acc_data_17_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_2, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1626_nl = MUX_s_1_2_2(buf_acc_data_17_17_0_sva,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign buf_acc_data_17_17_0_sva_dfm_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1626_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_1_slc_buf_acc_data_57_56_0_sat_sva_56_46_1
      = MUX_v_11_324_2(buf_acc_data_0_0_56_46_sva_dfm_1, buf_acc_data_0_1_56_46_sva_dfm_1,
      buf_acc_data_0_2_56_46_sva_dfm_1, buf_acc_data_0_3_56_46_sva_dfm_1, buf_acc_data_0_4_56_46_sva_dfm_1,
      buf_acc_data_0_5_56_46_sva_dfm_1, buf_acc_data_0_6_56_46_sva_dfm_1, buf_acc_data_0_7_56_46_sva_dfm_1,
      buf_acc_data_0_8_56_46_sva_dfm_1, buf_acc_data_0_9_56_46_sva_dfm_1, buf_acc_data_0_10_56_46_sva_dfm_1,
      buf_acc_data_0_11_56_46_sva_dfm_1, buf_acc_data_0_12_56_46_sva_dfm_1, buf_acc_data_0_13_56_46_sva_dfm_1,
      buf_acc_data_0_14_56_46_sva_dfm_1, buf_acc_data_0_15_56_46_sva_dfm_1, buf_acc_data_0_16_56_46_sva_dfm_1,
      buf_acc_data_0_17_56_46_sva_dfm_1, buf_acc_data_1_0_56_46_sva_dfm_1, buf_acc_data_1_1_56_46_sva_dfm_1,
      buf_acc_data_1_2_56_46_sva_dfm_1, buf_acc_data_1_3_56_46_sva_dfm_1, buf_acc_data_1_4_56_46_sva_dfm_1,
      buf_acc_data_1_5_56_46_sva_dfm_1, buf_acc_data_1_6_56_46_sva_dfm_1, buf_acc_data_1_7_56_46_sva_dfm_1,
      buf_acc_data_1_8_56_46_sva_dfm_1, buf_acc_data_1_9_56_46_sva_dfm_1, buf_acc_data_1_10_56_46_sva_dfm_1,
      buf_acc_data_1_11_56_46_sva_dfm_1, buf_acc_data_1_12_56_46_sva_dfm_1, buf_acc_data_1_13_56_46_sva_dfm_1,
      buf_acc_data_1_14_56_46_sva_dfm_1, buf_acc_data_1_15_56_46_sva_dfm_1, buf_acc_data_1_16_56_46_sva_dfm_1,
      buf_acc_data_1_17_56_46_sva_dfm_1, buf_acc_data_2_0_56_46_sva_dfm_1, buf_acc_data_2_1_56_46_sva_dfm_1,
      buf_acc_data_2_2_56_46_sva_dfm_1, buf_acc_data_2_3_56_46_sva_dfm_1, buf_acc_data_2_4_56_46_sva_dfm_1,
      buf_acc_data_2_5_56_46_sva_dfm_1, buf_acc_data_2_6_56_46_sva_dfm_1, buf_acc_data_2_7_56_46_sva_dfm_1,
      buf_acc_data_2_8_56_46_sva_dfm_1, buf_acc_data_2_9_56_46_sva_dfm_1, buf_acc_data_2_10_56_46_sva_dfm_1,
      buf_acc_data_2_11_56_46_sva_dfm_1, buf_acc_data_2_12_56_46_sva_dfm_1, buf_acc_data_2_13_56_46_sva_dfm_1,
      buf_acc_data_2_14_56_46_sva_dfm_1, buf_acc_data_2_15_56_46_sva_dfm_1, buf_acc_data_2_16_56_46_sva_dfm_1,
      buf_acc_data_2_17_56_46_sva_dfm_1, buf_acc_data_3_0_56_46_sva_dfm_1, buf_acc_data_3_1_56_46_sva_dfm_1,
      buf_acc_data_3_2_56_46_sva_dfm_1, buf_acc_data_3_3_56_46_sva_dfm_1, buf_acc_data_3_4_56_46_sva_dfm_1,
      buf_acc_data_3_5_56_46_sva_dfm_1, buf_acc_data_3_6_56_46_sva_dfm_1, buf_acc_data_3_7_56_46_sva_dfm_1,
      buf_acc_data_3_8_56_46_sva_dfm_1, buf_acc_data_3_9_56_46_sva_dfm_1, buf_acc_data_3_10_56_46_sva_dfm_1,
      buf_acc_data_3_11_56_46_sva_dfm_1, buf_acc_data_3_12_56_46_sva_dfm_1, buf_acc_data_3_13_56_46_sva_dfm_1,
      buf_acc_data_3_14_56_46_sva_dfm_1, buf_acc_data_3_15_56_46_sva_dfm_1, buf_acc_data_3_16_56_46_sva_dfm_1,
      buf_acc_data_3_17_56_46_sva_dfm_1, buf_acc_data_4_0_56_46_sva_dfm_1, buf_acc_data_4_1_56_46_sva_dfm_1,
      buf_acc_data_4_2_56_46_sva_dfm_1, buf_acc_data_4_3_56_46_sva_dfm_1, buf_acc_data_4_4_56_46_sva_dfm_1,
      buf_acc_data_4_5_56_46_sva_dfm_1, buf_acc_data_4_6_56_46_sva_dfm_1, buf_acc_data_4_7_56_46_sva_dfm_1,
      buf_acc_data_4_8_56_46_sva_dfm_1, buf_acc_data_4_9_56_46_sva_dfm_1, buf_acc_data_4_10_56_46_sva_dfm_1,
      buf_acc_data_4_11_56_46_sva_dfm_1, buf_acc_data_4_12_56_46_sva_dfm_1, buf_acc_data_4_13_56_46_sva_dfm_1,
      buf_acc_data_4_14_56_46_sva_dfm_1, buf_acc_data_4_15_56_46_sva_dfm_1, buf_acc_data_4_16_56_46_sva_dfm_1,
      buf_acc_data_4_17_56_46_sva_dfm_1, buf_acc_data_5_0_56_46_sva_dfm_1, buf_acc_data_5_1_56_46_sva_dfm_1,
      buf_acc_data_5_2_56_46_sva_dfm_1, buf_acc_data_5_3_56_46_sva_dfm_1, buf_acc_data_5_4_56_46_sva_dfm_1,
      buf_acc_data_5_5_56_46_sva_dfm_1, buf_acc_data_5_6_56_46_sva_dfm_1, buf_acc_data_5_7_56_46_sva_dfm_1,
      buf_acc_data_5_8_56_46_sva_dfm_1, buf_acc_data_5_9_56_46_sva_dfm_1, buf_acc_data_5_10_56_46_sva_dfm_1,
      buf_acc_data_5_11_56_46_sva_dfm_1, buf_acc_data_5_12_56_46_sva_dfm_1, buf_acc_data_5_13_56_46_sva_dfm_1,
      buf_acc_data_5_14_56_46_sva_dfm_1, buf_acc_data_5_15_56_46_sva_dfm_1, buf_acc_data_5_16_56_46_sva_dfm_1,
      buf_acc_data_5_17_56_46_sva_dfm_1, buf_acc_data_6_0_56_46_sva_dfm_1, buf_acc_data_6_1_56_46_sva_dfm_1,
      buf_acc_data_6_2_56_46_sva_dfm_1, buf_acc_data_6_3_56_46_sva_dfm_1, buf_acc_data_6_4_56_46_sva_dfm_1,
      buf_acc_data_6_5_56_46_sva_dfm_1, buf_acc_data_6_6_56_46_sva_dfm_1, buf_acc_data_6_7_56_46_sva_dfm_1,
      buf_acc_data_6_8_56_46_sva_dfm_1, buf_acc_data_6_9_56_46_sva_dfm_1, buf_acc_data_6_10_56_46_sva_dfm_1,
      buf_acc_data_6_11_56_46_sva_dfm_1, buf_acc_data_6_12_56_46_sva_dfm_1, buf_acc_data_6_13_56_46_sva_dfm_1,
      buf_acc_data_6_14_56_46_sva_dfm_1, buf_acc_data_6_15_56_46_sva_dfm_1, buf_acc_data_6_16_56_46_sva_dfm_1,
      buf_acc_data_6_17_56_46_sva_dfm_1, buf_acc_data_7_0_56_46_sva_dfm_1, buf_acc_data_7_1_56_46_sva_dfm_1,
      buf_acc_data_7_2_56_46_sva_dfm_1, buf_acc_data_7_3_56_46_sva_dfm_1, buf_acc_data_7_4_56_46_sva_dfm_1,
      buf_acc_data_7_5_56_46_sva_dfm_1, buf_acc_data_7_6_56_46_sva_dfm_1, buf_acc_data_7_7_56_46_sva_dfm_1,
      buf_acc_data_7_8_56_46_sva_dfm_1, buf_acc_data_7_9_56_46_sva_dfm_1, buf_acc_data_7_10_56_46_sva_dfm_1,
      buf_acc_data_7_11_56_46_sva_dfm_1, buf_acc_data_7_12_56_46_sva_dfm_1, buf_acc_data_7_13_56_46_sva_dfm_1,
      buf_acc_data_7_14_56_46_sva_dfm_1, buf_acc_data_7_15_56_46_sva_dfm_1, buf_acc_data_7_16_56_46_sva_dfm_1,
      buf_acc_data_7_17_56_46_sva_dfm_1, buf_acc_data_8_0_56_46_sva_dfm_1, buf_acc_data_8_1_56_46_sva_dfm_1,
      buf_acc_data_8_2_56_46_sva_dfm_1, buf_acc_data_8_3_56_46_sva_dfm_1, buf_acc_data_8_4_56_46_sva_dfm_1,
      buf_acc_data_8_5_56_46_sva_dfm_1, buf_acc_data_8_6_56_46_sva_dfm_1, buf_acc_data_8_7_56_46_sva_dfm_1,
      buf_acc_data_8_8_56_46_sva_dfm_1, buf_acc_data_8_9_56_46_sva_dfm_1, buf_acc_data_8_10_56_46_sva_dfm_1,
      buf_acc_data_8_11_56_46_sva_dfm_1, buf_acc_data_8_12_56_46_sva_dfm_1, buf_acc_data_8_13_56_46_sva_dfm_1,
      buf_acc_data_8_14_56_46_sva_dfm_1, buf_acc_data_8_15_56_46_sva_dfm_1, buf_acc_data_8_16_56_46_sva_dfm_1,
      buf_acc_data_8_17_56_46_sva_dfm_1, buf_acc_data_9_0_56_46_sva_dfm_1, buf_acc_data_9_1_56_46_sva_dfm_1,
      buf_acc_data_9_2_56_46_sva_dfm_1, buf_acc_data_9_3_56_46_sva_dfm_1, buf_acc_data_9_4_56_46_sva_dfm_1,
      buf_acc_data_9_5_56_46_sva_dfm_1, buf_acc_data_9_6_56_46_sva_dfm_1, buf_acc_data_9_7_56_46_sva_dfm_1,
      buf_acc_data_9_8_56_46_sva_dfm_1, buf_acc_data_9_9_56_46_sva_dfm_1, buf_acc_data_9_10_56_46_sva_dfm_1,
      buf_acc_data_9_11_56_46_sva_dfm_1, buf_acc_data_9_12_56_46_sva_dfm_1, buf_acc_data_9_13_56_46_sva_dfm_1,
      buf_acc_data_9_14_56_46_sva_dfm_1, buf_acc_data_9_15_56_46_sva_dfm_1, buf_acc_data_9_16_56_46_sva_dfm_1,
      buf_acc_data_9_17_56_46_sva_dfm_1, buf_acc_data_10_0_56_46_sva_dfm_1, buf_acc_data_10_1_56_46_sva_dfm_1,
      buf_acc_data_10_2_56_46_sva_dfm_1, buf_acc_data_10_3_56_46_sva_dfm_1, buf_acc_data_10_4_56_46_sva_dfm_1,
      buf_acc_data_10_5_56_46_sva_dfm_1, buf_acc_data_10_6_56_46_sva_dfm_1, buf_acc_data_10_7_56_46_sva_dfm_1,
      buf_acc_data_10_8_56_46_sva_dfm_1, buf_acc_data_10_9_56_46_sva_dfm_1, buf_acc_data_10_10_56_46_sva_dfm_1,
      buf_acc_data_10_11_56_46_sva_dfm_1, buf_acc_data_10_12_56_46_sva_dfm_1, buf_acc_data_10_13_56_46_sva_dfm_1,
      buf_acc_data_10_14_56_46_sva_dfm_1, buf_acc_data_10_15_56_46_sva_dfm_1, buf_acc_data_10_16_56_46_sva_dfm_1,
      buf_acc_data_10_17_56_46_sva_dfm_1, buf_acc_data_11_0_56_46_sva_dfm_1, buf_acc_data_11_1_56_46_sva_dfm_1,
      buf_acc_data_11_2_56_46_sva_dfm_1, buf_acc_data_11_3_56_46_sva_dfm_1, buf_acc_data_11_4_56_46_sva_dfm_1,
      buf_acc_data_11_5_56_46_sva_dfm_1, buf_acc_data_11_6_56_46_sva_dfm_1, buf_acc_data_11_7_56_46_sva_dfm_1,
      buf_acc_data_11_8_56_46_sva_dfm_1, buf_acc_data_11_9_56_46_sva_dfm_1, buf_acc_data_11_10_56_46_sva_dfm_1,
      buf_acc_data_11_11_56_46_sva_dfm_1, buf_acc_data_11_12_56_46_sva_dfm_1, buf_acc_data_11_13_56_46_sva_dfm_1,
      buf_acc_data_11_14_56_46_sva_dfm_1, buf_acc_data_11_15_56_46_sva_dfm_1, buf_acc_data_11_16_56_46_sva_dfm_1,
      buf_acc_data_11_17_56_46_sva_dfm_1, buf_acc_data_12_0_56_46_sva_dfm_1, buf_acc_data_12_1_56_46_sva_dfm_1,
      buf_acc_data_12_2_56_46_sva_dfm_1, buf_acc_data_12_3_56_46_sva_dfm_1, buf_acc_data_12_4_56_46_sva_dfm_1,
      buf_acc_data_12_5_56_46_sva_dfm_1, buf_acc_data_12_6_56_46_sva_dfm_1, buf_acc_data_12_7_56_46_sva_dfm_1,
      buf_acc_data_12_8_56_46_sva_dfm_1, buf_acc_data_12_9_56_46_sva_dfm_1, buf_acc_data_12_10_56_46_sva_dfm_1,
      buf_acc_data_12_11_56_46_sva_dfm_1, buf_acc_data_12_12_56_46_sva_dfm_1, buf_acc_data_12_13_56_46_sva_dfm_1,
      buf_acc_data_12_14_56_46_sva_dfm_1, buf_acc_data_12_15_56_46_sva_dfm_1, buf_acc_data_12_16_56_46_sva_dfm_1,
      buf_acc_data_12_17_56_46_sva_dfm_1, buf_acc_data_13_0_56_46_sva_dfm_1, buf_acc_data_13_1_56_46_sva_dfm_1,
      buf_acc_data_13_2_56_46_sva_dfm_1, buf_acc_data_13_3_56_46_sva_dfm_1, buf_acc_data_13_4_56_46_sva_dfm_1,
      buf_acc_data_13_5_56_46_sva_dfm_1, buf_acc_data_13_6_56_46_sva_dfm_1, buf_acc_data_13_7_56_46_sva_dfm_1,
      buf_acc_data_13_8_56_46_sva_dfm_1, buf_acc_data_13_9_56_46_sva_dfm_1, buf_acc_data_13_10_56_46_sva_dfm_1,
      buf_acc_data_13_11_56_46_sva_dfm_1, buf_acc_data_13_12_56_46_sva_dfm_1, buf_acc_data_13_13_56_46_sva_dfm_1,
      buf_acc_data_13_14_56_46_sva_dfm_1, buf_acc_data_13_15_56_46_sva_dfm_1, buf_acc_data_13_16_56_46_sva_dfm_1,
      buf_acc_data_13_17_56_46_sva_dfm_1, buf_acc_data_14_0_56_46_sva_dfm_1, buf_acc_data_14_1_56_46_sva_dfm_1,
      buf_acc_data_14_2_56_46_sva_dfm_1, buf_acc_data_14_3_56_46_sva_dfm_1, buf_acc_data_14_4_56_46_sva_dfm_1,
      buf_acc_data_14_5_56_46_sva_dfm_1, buf_acc_data_14_6_56_46_sva_dfm_1, buf_acc_data_14_7_56_46_sva_dfm_1,
      buf_acc_data_14_8_56_46_sva_dfm_1, buf_acc_data_14_9_56_46_sva_dfm_1, buf_acc_data_14_10_56_46_sva_dfm_1,
      buf_acc_data_14_11_56_46_sva_dfm_1, buf_acc_data_14_12_56_46_sva_dfm_1, buf_acc_data_14_13_56_46_sva_dfm_1,
      buf_acc_data_14_14_56_46_sva_dfm_1, buf_acc_data_14_15_56_46_sva_dfm_1, buf_acc_data_14_16_56_46_sva_dfm_1,
      buf_acc_data_14_17_56_46_sva_dfm_1, buf_acc_data_15_0_56_46_sva_dfm_1, buf_acc_data_15_1_56_46_sva_dfm_1,
      buf_acc_data_15_2_56_46_sva_dfm_1, buf_acc_data_15_3_56_46_sva_dfm_1, buf_acc_data_15_4_56_46_sva_dfm_1,
      buf_acc_data_15_5_56_46_sva_dfm_1, buf_acc_data_15_6_56_46_sva_dfm_1, buf_acc_data_15_7_56_46_sva_dfm_1,
      buf_acc_data_15_8_56_46_sva_dfm_1, buf_acc_data_15_9_56_46_sva_dfm_1, buf_acc_data_15_10_56_46_sva_dfm_1,
      buf_acc_data_15_11_56_46_sva_dfm_1, buf_acc_data_15_12_56_46_sva_dfm_1, buf_acc_data_15_13_56_46_sva_dfm_1,
      buf_acc_data_15_14_56_46_sva_dfm_1, buf_acc_data_15_15_56_46_sva_dfm_1, buf_acc_data_15_16_56_46_sva_dfm_1,
      buf_acc_data_15_17_56_46_sva_dfm_1, buf_acc_data_16_0_56_46_sva_dfm_1, buf_acc_data_16_1_56_46_sva_dfm_1,
      buf_acc_data_16_2_56_46_sva_dfm_1, buf_acc_data_16_3_56_46_sva_dfm_1, buf_acc_data_16_4_56_46_sva_dfm_1,
      buf_acc_data_16_5_56_46_sva_dfm_1, buf_acc_data_16_6_56_46_sva_dfm_1, buf_acc_data_16_7_56_46_sva_dfm_1,
      buf_acc_data_16_8_56_46_sva_dfm_1, buf_acc_data_16_9_56_46_sva_dfm_1, buf_acc_data_16_10_56_46_sva_dfm_1,
      buf_acc_data_16_11_56_46_sva_dfm_1, buf_acc_data_16_12_56_46_sva_dfm_1, buf_acc_data_16_13_56_46_sva_dfm_1,
      buf_acc_data_16_14_56_46_sva_dfm_1, buf_acc_data_16_15_56_46_sva_dfm_1, buf_acc_data_16_16_56_46_sva_dfm_1,
      buf_acc_data_16_17_56_46_sva_dfm_1, buf_acc_data_17_0_56_46_sva_dfm_1, buf_acc_data_17_1_56_46_sva_dfm_1,
      buf_acc_data_17_2_56_46_sva_dfm_1, buf_acc_data_17_3_56_46_sva_dfm_1, buf_acc_data_17_4_56_46_sva_dfm_1,
      buf_acc_data_17_5_56_46_sva_dfm_1, buf_acc_data_17_6_56_46_sva_dfm_1, buf_acc_data_17_7_56_46_sva_dfm_1,
      buf_acc_data_17_8_56_46_sva_dfm_1, buf_acc_data_17_9_56_46_sva_dfm_1, buf_acc_data_17_10_56_46_sva_dfm_1,
      buf_acc_data_17_11_56_46_sva_dfm_1, buf_acc_data_17_12_56_46_sva_dfm_1, buf_acc_data_17_13_56_46_sva_dfm_1,
      buf_acc_data_17_14_56_46_sva_dfm_1, buf_acc_data_17_15_56_46_sva_dfm_1, buf_acc_data_17_16_56_46_sva_dfm_1,
      buf_acc_data_17_17_56_46_sva_dfm_1, {CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_2
      , CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_2
      , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0});
  assign buf_acc_data_0_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5508
      , CONVOLUTION_LOOP_for_for_for_asn_5510 , CONVOLUTION_LOOP_for_for_for_asn_5512});
  assign buf_acc_data_0_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5502
      , CONVOLUTION_LOOP_for_for_for_asn_5504 , CONVOLUTION_LOOP_for_for_for_asn_5506});
  assign buf_acc_data_0_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5496
      , CONVOLUTION_LOOP_for_for_for_asn_5498 , CONVOLUTION_LOOP_for_for_for_asn_5500});
  assign buf_acc_data_0_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5490
      , CONVOLUTION_LOOP_for_for_for_asn_5492 , CONVOLUTION_LOOP_for_for_for_asn_5494});
  assign buf_acc_data_0_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5484
      , CONVOLUTION_LOOP_for_for_for_asn_5486 , CONVOLUTION_LOOP_for_for_for_asn_5488});
  assign buf_acc_data_0_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5478
      , CONVOLUTION_LOOP_for_for_for_asn_5480 , CONVOLUTION_LOOP_for_for_for_asn_5482});
  assign buf_acc_data_0_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5472
      , CONVOLUTION_LOOP_for_for_for_asn_5474 , CONVOLUTION_LOOP_for_for_for_asn_5476});
  assign buf_acc_data_0_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5466
      , CONVOLUTION_LOOP_for_for_for_asn_5468 , CONVOLUTION_LOOP_for_for_for_asn_5470});
  assign buf_acc_data_0_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5460
      , CONVOLUTION_LOOP_for_for_for_asn_5462 , CONVOLUTION_LOOP_for_for_for_asn_5464});
  assign buf_acc_data_0_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5454
      , CONVOLUTION_LOOP_for_for_for_asn_5456 , CONVOLUTION_LOOP_for_for_for_asn_5458});
  assign buf_acc_data_0_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5448
      , CONVOLUTION_LOOP_for_for_for_asn_5450 , CONVOLUTION_LOOP_for_for_for_asn_5452});
  assign buf_acc_data_0_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5442
      , CONVOLUTION_LOOP_for_for_for_asn_5444 , CONVOLUTION_LOOP_for_for_for_asn_5446});
  assign buf_acc_data_0_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5436
      , CONVOLUTION_LOOP_for_for_for_asn_5438 , CONVOLUTION_LOOP_for_for_for_asn_5440});
  assign buf_acc_data_0_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5430
      , CONVOLUTION_LOOP_for_for_for_asn_5432 , CONVOLUTION_LOOP_for_for_for_asn_5434});
  assign buf_acc_data_0_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5424
      , CONVOLUTION_LOOP_for_for_for_asn_5426 , CONVOLUTION_LOOP_for_for_for_asn_5428});
  assign buf_acc_data_0_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5418
      , CONVOLUTION_LOOP_for_for_for_asn_5420 , CONVOLUTION_LOOP_for_for_for_asn_5422});
  assign buf_acc_data_0_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5412
      , CONVOLUTION_LOOP_for_for_for_asn_5414 , CONVOLUTION_LOOP_for_for_for_asn_5416});
  assign buf_acc_data_0_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_0_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5406
      , CONVOLUTION_LOOP_for_for_for_asn_5408 , CONVOLUTION_LOOP_for_for_for_asn_5410});
  assign buf_acc_data_1_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5400
      , CONVOLUTION_LOOP_for_for_for_asn_5402 , CONVOLUTION_LOOP_for_for_for_asn_5404});
  assign buf_acc_data_1_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5394
      , CONVOLUTION_LOOP_for_for_for_asn_5396 , CONVOLUTION_LOOP_for_for_for_asn_5398});
  assign buf_acc_data_1_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5388
      , CONVOLUTION_LOOP_for_for_for_asn_5390 , CONVOLUTION_LOOP_for_for_for_asn_5392});
  assign buf_acc_data_1_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5382
      , CONVOLUTION_LOOP_for_for_for_asn_5384 , CONVOLUTION_LOOP_for_for_for_asn_5386});
  assign buf_acc_data_1_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5376
      , CONVOLUTION_LOOP_for_for_for_asn_5378 , CONVOLUTION_LOOP_for_for_for_asn_5380});
  assign buf_acc_data_1_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5370
      , CONVOLUTION_LOOP_for_for_for_asn_5372 , CONVOLUTION_LOOP_for_for_for_asn_5374});
  assign buf_acc_data_1_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5364
      , CONVOLUTION_LOOP_for_for_for_asn_5366 , CONVOLUTION_LOOP_for_for_for_asn_5368});
  assign buf_acc_data_1_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5358
      , CONVOLUTION_LOOP_for_for_for_asn_5360 , CONVOLUTION_LOOP_for_for_for_asn_5362});
  assign buf_acc_data_1_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5352
      , CONVOLUTION_LOOP_for_for_for_asn_5354 , CONVOLUTION_LOOP_for_for_for_asn_5356});
  assign buf_acc_data_1_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5346
      , CONVOLUTION_LOOP_for_for_for_asn_5348 , CONVOLUTION_LOOP_for_for_for_asn_5350});
  assign buf_acc_data_1_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5340
      , CONVOLUTION_LOOP_for_for_for_asn_5342 , CONVOLUTION_LOOP_for_for_for_asn_5344});
  assign buf_acc_data_1_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5334
      , CONVOLUTION_LOOP_for_for_for_asn_5336 , CONVOLUTION_LOOP_for_for_for_asn_5338});
  assign buf_acc_data_1_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5328
      , CONVOLUTION_LOOP_for_for_for_asn_5330 , CONVOLUTION_LOOP_for_for_for_asn_5332});
  assign buf_acc_data_1_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5322
      , CONVOLUTION_LOOP_for_for_for_asn_5324 , CONVOLUTION_LOOP_for_for_for_asn_5326});
  assign buf_acc_data_1_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5316
      , CONVOLUTION_LOOP_for_for_for_asn_5318 , CONVOLUTION_LOOP_for_for_for_asn_5320});
  assign buf_acc_data_1_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5310
      , CONVOLUTION_LOOP_for_for_for_asn_5312 , CONVOLUTION_LOOP_for_for_for_asn_5314});
  assign buf_acc_data_1_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5304
      , CONVOLUTION_LOOP_for_for_for_asn_5306 , CONVOLUTION_LOOP_for_for_for_asn_5308});
  assign buf_acc_data_1_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_1_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5298
      , CONVOLUTION_LOOP_for_for_for_asn_5300 , CONVOLUTION_LOOP_for_for_for_asn_5302});
  assign buf_acc_data_2_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5292
      , CONVOLUTION_LOOP_for_for_for_asn_5294 , CONVOLUTION_LOOP_for_for_for_asn_5296});
  assign buf_acc_data_2_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5286
      , CONVOLUTION_LOOP_for_for_for_asn_5288 , CONVOLUTION_LOOP_for_for_for_asn_5290});
  assign buf_acc_data_2_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5280
      , CONVOLUTION_LOOP_for_for_for_asn_5282 , CONVOLUTION_LOOP_for_for_for_asn_5284});
  assign buf_acc_data_2_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5274
      , CONVOLUTION_LOOP_for_for_for_asn_5276 , CONVOLUTION_LOOP_for_for_for_asn_5278});
  assign buf_acc_data_2_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5268
      , CONVOLUTION_LOOP_for_for_for_asn_5270 , CONVOLUTION_LOOP_for_for_for_asn_5272});
  assign buf_acc_data_2_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5262
      , CONVOLUTION_LOOP_for_for_for_asn_5264 , CONVOLUTION_LOOP_for_for_for_asn_5266});
  assign buf_acc_data_2_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5256
      , CONVOLUTION_LOOP_for_for_for_asn_5258 , CONVOLUTION_LOOP_for_for_for_asn_5260});
  assign buf_acc_data_2_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5250
      , CONVOLUTION_LOOP_for_for_for_asn_5252 , CONVOLUTION_LOOP_for_for_for_asn_5254});
  assign buf_acc_data_2_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5244
      , CONVOLUTION_LOOP_for_for_for_asn_5246 , CONVOLUTION_LOOP_for_for_for_asn_5248});
  assign buf_acc_data_2_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5238
      , CONVOLUTION_LOOP_for_for_for_asn_5240 , CONVOLUTION_LOOP_for_for_for_asn_5242});
  assign buf_acc_data_2_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5232
      , CONVOLUTION_LOOP_for_for_for_asn_5234 , CONVOLUTION_LOOP_for_for_for_asn_5236});
  assign buf_acc_data_2_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5226
      , CONVOLUTION_LOOP_for_for_for_asn_5228 , CONVOLUTION_LOOP_for_for_for_asn_5230});
  assign buf_acc_data_2_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5220
      , CONVOLUTION_LOOP_for_for_for_asn_5222 , CONVOLUTION_LOOP_for_for_for_asn_5224});
  assign buf_acc_data_2_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5214
      , CONVOLUTION_LOOP_for_for_for_asn_5216 , CONVOLUTION_LOOP_for_for_for_asn_5218});
  assign buf_acc_data_2_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5208
      , CONVOLUTION_LOOP_for_for_for_asn_5210 , CONVOLUTION_LOOP_for_for_for_asn_5212});
  assign buf_acc_data_2_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5202
      , CONVOLUTION_LOOP_for_for_for_asn_5204 , CONVOLUTION_LOOP_for_for_for_asn_5206});
  assign buf_acc_data_2_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5196
      , CONVOLUTION_LOOP_for_for_for_asn_5198 , CONVOLUTION_LOOP_for_for_for_asn_5200});
  assign buf_acc_data_2_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_2_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5190
      , CONVOLUTION_LOOP_for_for_for_asn_5192 , CONVOLUTION_LOOP_for_for_for_asn_5194});
  assign buf_acc_data_3_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5184
      , CONVOLUTION_LOOP_for_for_for_asn_5186 , CONVOLUTION_LOOP_for_for_for_asn_5188});
  assign buf_acc_data_3_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5178
      , CONVOLUTION_LOOP_for_for_for_asn_5180 , CONVOLUTION_LOOP_for_for_for_asn_5182});
  assign buf_acc_data_3_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5172
      , CONVOLUTION_LOOP_for_for_for_asn_5174 , CONVOLUTION_LOOP_for_for_for_asn_5176});
  assign buf_acc_data_3_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5166
      , CONVOLUTION_LOOP_for_for_for_asn_5168 , CONVOLUTION_LOOP_for_for_for_asn_5170});
  assign buf_acc_data_3_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5160
      , CONVOLUTION_LOOP_for_for_for_asn_5162 , CONVOLUTION_LOOP_for_for_for_asn_5164});
  assign buf_acc_data_3_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5154
      , CONVOLUTION_LOOP_for_for_for_asn_5156 , CONVOLUTION_LOOP_for_for_for_asn_5158});
  assign buf_acc_data_3_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5148
      , CONVOLUTION_LOOP_for_for_for_asn_5150 , CONVOLUTION_LOOP_for_for_for_asn_5152});
  assign buf_acc_data_3_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5142
      , CONVOLUTION_LOOP_for_for_for_asn_5144 , CONVOLUTION_LOOP_for_for_for_asn_5146});
  assign buf_acc_data_3_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5136
      , CONVOLUTION_LOOP_for_for_for_asn_5138 , CONVOLUTION_LOOP_for_for_for_asn_5140});
  assign buf_acc_data_3_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5130
      , CONVOLUTION_LOOP_for_for_for_asn_5132 , CONVOLUTION_LOOP_for_for_for_asn_5134});
  assign buf_acc_data_3_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5124
      , CONVOLUTION_LOOP_for_for_for_asn_5126 , CONVOLUTION_LOOP_for_for_for_asn_5128});
  assign buf_acc_data_3_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5118
      , CONVOLUTION_LOOP_for_for_for_asn_5120 , CONVOLUTION_LOOP_for_for_for_asn_5122});
  assign buf_acc_data_3_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5112
      , CONVOLUTION_LOOP_for_for_for_asn_5114 , CONVOLUTION_LOOP_for_for_for_asn_5116});
  assign buf_acc_data_3_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5106
      , CONVOLUTION_LOOP_for_for_for_asn_5108 , CONVOLUTION_LOOP_for_for_for_asn_5110});
  assign buf_acc_data_3_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5100
      , CONVOLUTION_LOOP_for_for_for_asn_5102 , CONVOLUTION_LOOP_for_for_for_asn_5104});
  assign buf_acc_data_3_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5094
      , CONVOLUTION_LOOP_for_for_for_asn_5096 , CONVOLUTION_LOOP_for_for_for_asn_5098});
  assign buf_acc_data_3_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5088
      , CONVOLUTION_LOOP_for_for_for_asn_5090 , CONVOLUTION_LOOP_for_for_for_asn_5092});
  assign buf_acc_data_3_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_3_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5082
      , CONVOLUTION_LOOP_for_for_for_asn_5084 , CONVOLUTION_LOOP_for_for_for_asn_5086});
  assign buf_acc_data_4_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5076
      , CONVOLUTION_LOOP_for_for_for_asn_5078 , CONVOLUTION_LOOP_for_for_for_asn_5080});
  assign buf_acc_data_4_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5070
      , CONVOLUTION_LOOP_for_for_for_asn_5072 , CONVOLUTION_LOOP_for_for_for_asn_5074});
  assign buf_acc_data_4_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5064
      , CONVOLUTION_LOOP_for_for_for_asn_5066 , CONVOLUTION_LOOP_for_for_for_asn_5068});
  assign buf_acc_data_4_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5058
      , CONVOLUTION_LOOP_for_for_for_asn_5060 , CONVOLUTION_LOOP_for_for_for_asn_5062});
  assign buf_acc_data_4_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5052
      , CONVOLUTION_LOOP_for_for_for_asn_5054 , CONVOLUTION_LOOP_for_for_for_asn_5056});
  assign buf_acc_data_4_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5046
      , CONVOLUTION_LOOP_for_for_for_asn_5048 , CONVOLUTION_LOOP_for_for_for_asn_5050});
  assign buf_acc_data_4_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5040
      , CONVOLUTION_LOOP_for_for_for_asn_5042 , CONVOLUTION_LOOP_for_for_for_asn_5044});
  assign buf_acc_data_4_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5034
      , CONVOLUTION_LOOP_for_for_for_asn_5036 , CONVOLUTION_LOOP_for_for_for_asn_5038});
  assign buf_acc_data_4_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5028
      , CONVOLUTION_LOOP_for_for_for_asn_5030 , CONVOLUTION_LOOP_for_for_for_asn_5032});
  assign buf_acc_data_4_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5022
      , CONVOLUTION_LOOP_for_for_for_asn_5024 , CONVOLUTION_LOOP_for_for_for_asn_5026});
  assign buf_acc_data_4_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5016
      , CONVOLUTION_LOOP_for_for_for_asn_5018 , CONVOLUTION_LOOP_for_for_for_asn_5020});
  assign buf_acc_data_4_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5010
      , CONVOLUTION_LOOP_for_for_for_asn_5012 , CONVOLUTION_LOOP_for_for_for_asn_5014});
  assign buf_acc_data_4_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5004
      , CONVOLUTION_LOOP_for_for_for_asn_5006 , CONVOLUTION_LOOP_for_for_for_asn_5008});
  assign buf_acc_data_4_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4998
      , CONVOLUTION_LOOP_for_for_for_asn_5000 , CONVOLUTION_LOOP_for_for_for_asn_5002});
  assign buf_acc_data_4_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4992
      , CONVOLUTION_LOOP_for_for_for_asn_4994 , CONVOLUTION_LOOP_for_for_for_asn_4996});
  assign buf_acc_data_4_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4986
      , CONVOLUTION_LOOP_for_for_for_asn_4988 , CONVOLUTION_LOOP_for_for_for_asn_4990});
  assign buf_acc_data_4_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4980
      , CONVOLUTION_LOOP_for_for_for_asn_4982 , CONVOLUTION_LOOP_for_for_for_asn_4984});
  assign buf_acc_data_4_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_4_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4974
      , CONVOLUTION_LOOP_for_for_for_asn_4976 , CONVOLUTION_LOOP_for_for_for_asn_4978});
  assign buf_acc_data_5_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4968
      , CONVOLUTION_LOOP_for_for_for_asn_4970 , CONVOLUTION_LOOP_for_for_for_asn_4972});
  assign buf_acc_data_5_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4962
      , CONVOLUTION_LOOP_for_for_for_asn_4964 , CONVOLUTION_LOOP_for_for_for_asn_4966});
  assign buf_acc_data_5_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4956
      , CONVOLUTION_LOOP_for_for_for_asn_4958 , CONVOLUTION_LOOP_for_for_for_asn_4960});
  assign buf_acc_data_5_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4950
      , CONVOLUTION_LOOP_for_for_for_asn_4952 , CONVOLUTION_LOOP_for_for_for_asn_4954});
  assign buf_acc_data_5_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4944
      , CONVOLUTION_LOOP_for_for_for_asn_4946 , CONVOLUTION_LOOP_for_for_for_asn_4948});
  assign buf_acc_data_5_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4938
      , CONVOLUTION_LOOP_for_for_for_asn_4940 , CONVOLUTION_LOOP_for_for_for_asn_4942});
  assign buf_acc_data_5_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4932
      , CONVOLUTION_LOOP_for_for_for_asn_4934 , CONVOLUTION_LOOP_for_for_for_asn_4936});
  assign buf_acc_data_5_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4926
      , CONVOLUTION_LOOP_for_for_for_asn_4928 , CONVOLUTION_LOOP_for_for_for_asn_4930});
  assign buf_acc_data_5_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4920
      , CONVOLUTION_LOOP_for_for_for_asn_4922 , CONVOLUTION_LOOP_for_for_for_asn_4924});
  assign buf_acc_data_5_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4914
      , CONVOLUTION_LOOP_for_for_for_asn_4916 , CONVOLUTION_LOOP_for_for_for_asn_4918});
  assign buf_acc_data_5_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4908
      , CONVOLUTION_LOOP_for_for_for_asn_4910 , CONVOLUTION_LOOP_for_for_for_asn_4912});
  assign buf_acc_data_5_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4902
      , CONVOLUTION_LOOP_for_for_for_asn_4904 , CONVOLUTION_LOOP_for_for_for_asn_4906});
  assign buf_acc_data_5_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4896
      , CONVOLUTION_LOOP_for_for_for_asn_4898 , CONVOLUTION_LOOP_for_for_for_asn_4900});
  assign buf_acc_data_5_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4890
      , CONVOLUTION_LOOP_for_for_for_asn_4892 , CONVOLUTION_LOOP_for_for_for_asn_4894});
  assign buf_acc_data_5_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4884
      , CONVOLUTION_LOOP_for_for_for_asn_4886 , CONVOLUTION_LOOP_for_for_for_asn_4888});
  assign buf_acc_data_5_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4878
      , CONVOLUTION_LOOP_for_for_for_asn_4880 , CONVOLUTION_LOOP_for_for_for_asn_4882});
  assign buf_acc_data_5_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4872
      , CONVOLUTION_LOOP_for_for_for_asn_4874 , CONVOLUTION_LOOP_for_for_for_asn_4876});
  assign buf_acc_data_5_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_5_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4866
      , CONVOLUTION_LOOP_for_for_for_asn_4868 , CONVOLUTION_LOOP_for_for_for_asn_4870});
  assign buf_acc_data_6_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4860
      , CONVOLUTION_LOOP_for_for_for_asn_4862 , CONVOLUTION_LOOP_for_for_for_asn_4864});
  assign buf_acc_data_6_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4854
      , CONVOLUTION_LOOP_for_for_for_asn_4856 , CONVOLUTION_LOOP_for_for_for_asn_4858});
  assign buf_acc_data_6_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4848
      , CONVOLUTION_LOOP_for_for_for_asn_4850 , CONVOLUTION_LOOP_for_for_for_asn_4852});
  assign buf_acc_data_6_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4842
      , CONVOLUTION_LOOP_for_for_for_asn_4844 , CONVOLUTION_LOOP_for_for_for_asn_4846});
  assign buf_acc_data_6_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4836
      , CONVOLUTION_LOOP_for_for_for_asn_4838 , CONVOLUTION_LOOP_for_for_for_asn_4840});
  assign buf_acc_data_6_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4830
      , CONVOLUTION_LOOP_for_for_for_asn_4832 , CONVOLUTION_LOOP_for_for_for_asn_4834});
  assign buf_acc_data_6_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4824
      , CONVOLUTION_LOOP_for_for_for_asn_4826 , CONVOLUTION_LOOP_for_for_for_asn_4828});
  assign buf_acc_data_6_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4818
      , CONVOLUTION_LOOP_for_for_for_asn_4820 , CONVOLUTION_LOOP_for_for_for_asn_4822});
  assign buf_acc_data_6_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4812
      , CONVOLUTION_LOOP_for_for_for_asn_4814 , CONVOLUTION_LOOP_for_for_for_asn_4816});
  assign buf_acc_data_6_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4806
      , CONVOLUTION_LOOP_for_for_for_asn_4808 , CONVOLUTION_LOOP_for_for_for_asn_4810});
  assign buf_acc_data_6_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4800
      , CONVOLUTION_LOOP_for_for_for_asn_4802 , CONVOLUTION_LOOP_for_for_for_asn_4804});
  assign buf_acc_data_6_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4794
      , CONVOLUTION_LOOP_for_for_for_asn_4796 , CONVOLUTION_LOOP_for_for_for_asn_4798});
  assign buf_acc_data_6_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4788
      , CONVOLUTION_LOOP_for_for_for_asn_4790 , CONVOLUTION_LOOP_for_for_for_asn_4792});
  assign buf_acc_data_6_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4782
      , CONVOLUTION_LOOP_for_for_for_asn_4784 , CONVOLUTION_LOOP_for_for_for_asn_4786});
  assign buf_acc_data_6_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4776
      , CONVOLUTION_LOOP_for_for_for_asn_4778 , CONVOLUTION_LOOP_for_for_for_asn_4780});
  assign buf_acc_data_6_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4770
      , CONVOLUTION_LOOP_for_for_for_asn_4772 , CONVOLUTION_LOOP_for_for_for_asn_4774});
  assign buf_acc_data_6_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4764
      , CONVOLUTION_LOOP_for_for_for_asn_4766 , CONVOLUTION_LOOP_for_for_for_asn_4768});
  assign buf_acc_data_6_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_6_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4758
      , CONVOLUTION_LOOP_for_for_for_asn_4760 , CONVOLUTION_LOOP_for_for_for_asn_4762});
  assign buf_acc_data_7_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4752
      , CONVOLUTION_LOOP_for_for_for_asn_4754 , CONVOLUTION_LOOP_for_for_for_asn_4756});
  assign buf_acc_data_7_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4746
      , CONVOLUTION_LOOP_for_for_for_asn_4748 , CONVOLUTION_LOOP_for_for_for_asn_4750});
  assign buf_acc_data_7_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4740
      , CONVOLUTION_LOOP_for_for_for_asn_4742 , CONVOLUTION_LOOP_for_for_for_asn_4744});
  assign buf_acc_data_7_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4734
      , CONVOLUTION_LOOP_for_for_for_asn_4736 , CONVOLUTION_LOOP_for_for_for_asn_4738});
  assign buf_acc_data_7_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4728
      , CONVOLUTION_LOOP_for_for_for_asn_4730 , CONVOLUTION_LOOP_for_for_for_asn_4732});
  assign buf_acc_data_7_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4722
      , CONVOLUTION_LOOP_for_for_for_asn_4724 , CONVOLUTION_LOOP_for_for_for_asn_4726});
  assign buf_acc_data_7_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4716
      , CONVOLUTION_LOOP_for_for_for_asn_4718 , CONVOLUTION_LOOP_for_for_for_asn_4720});
  assign buf_acc_data_7_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4710
      , CONVOLUTION_LOOP_for_for_for_asn_4712 , CONVOLUTION_LOOP_for_for_for_asn_4714});
  assign buf_acc_data_7_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4704
      , CONVOLUTION_LOOP_for_for_for_asn_4706 , CONVOLUTION_LOOP_for_for_for_asn_4708});
  assign buf_acc_data_7_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4698
      , CONVOLUTION_LOOP_for_for_for_asn_4700 , CONVOLUTION_LOOP_for_for_for_asn_4702});
  assign buf_acc_data_7_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4692
      , CONVOLUTION_LOOP_for_for_for_asn_4694 , CONVOLUTION_LOOP_for_for_for_asn_4696});
  assign buf_acc_data_7_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4686
      , CONVOLUTION_LOOP_for_for_for_asn_4688 , CONVOLUTION_LOOP_for_for_for_asn_4690});
  assign buf_acc_data_7_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4680
      , CONVOLUTION_LOOP_for_for_for_asn_4682 , CONVOLUTION_LOOP_for_for_for_asn_4684});
  assign buf_acc_data_7_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4674
      , CONVOLUTION_LOOP_for_for_for_asn_4676 , CONVOLUTION_LOOP_for_for_for_asn_4678});
  assign buf_acc_data_7_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4668
      , CONVOLUTION_LOOP_for_for_for_asn_4670 , CONVOLUTION_LOOP_for_for_for_asn_4672});
  assign buf_acc_data_7_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4662
      , CONVOLUTION_LOOP_for_for_for_asn_4664 , CONVOLUTION_LOOP_for_for_for_asn_4666});
  assign buf_acc_data_7_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4656
      , CONVOLUTION_LOOP_for_for_for_asn_4658 , CONVOLUTION_LOOP_for_for_for_asn_4660});
  assign buf_acc_data_7_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_7_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4650
      , CONVOLUTION_LOOP_for_for_for_asn_4652 , CONVOLUTION_LOOP_for_for_for_asn_4654});
  assign buf_acc_data_8_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4644
      , CONVOLUTION_LOOP_for_for_for_asn_4646 , CONVOLUTION_LOOP_for_for_for_asn_4648});
  assign buf_acc_data_8_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4638
      , CONVOLUTION_LOOP_for_for_for_asn_4640 , CONVOLUTION_LOOP_for_for_for_asn_4642});
  assign buf_acc_data_8_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4632
      , CONVOLUTION_LOOP_for_for_for_asn_4634 , CONVOLUTION_LOOP_for_for_for_asn_4636});
  assign buf_acc_data_8_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4626
      , CONVOLUTION_LOOP_for_for_for_asn_4628 , CONVOLUTION_LOOP_for_for_for_asn_4630});
  assign buf_acc_data_8_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4620
      , CONVOLUTION_LOOP_for_for_for_asn_4622 , CONVOLUTION_LOOP_for_for_for_asn_4624});
  assign buf_acc_data_8_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4614
      , CONVOLUTION_LOOP_for_for_for_asn_4616 , CONVOLUTION_LOOP_for_for_for_asn_4618});
  assign buf_acc_data_8_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4608
      , CONVOLUTION_LOOP_for_for_for_asn_4610 , CONVOLUTION_LOOP_for_for_for_asn_4612});
  assign buf_acc_data_8_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4602
      , CONVOLUTION_LOOP_for_for_for_asn_4604 , CONVOLUTION_LOOP_for_for_for_asn_4606});
  assign buf_acc_data_8_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4596
      , CONVOLUTION_LOOP_for_for_for_asn_4598 , CONVOLUTION_LOOP_for_for_for_asn_4600});
  assign buf_acc_data_8_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4590
      , CONVOLUTION_LOOP_for_for_for_asn_4592 , CONVOLUTION_LOOP_for_for_for_asn_4594});
  assign buf_acc_data_8_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4584
      , CONVOLUTION_LOOP_for_for_for_asn_4586 , CONVOLUTION_LOOP_for_for_for_asn_4588});
  assign buf_acc_data_8_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4578
      , CONVOLUTION_LOOP_for_for_for_asn_4580 , CONVOLUTION_LOOP_for_for_for_asn_4582});
  assign buf_acc_data_8_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4572
      , CONVOLUTION_LOOP_for_for_for_asn_4574 , CONVOLUTION_LOOP_for_for_for_asn_4576});
  assign buf_acc_data_8_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4566
      , CONVOLUTION_LOOP_for_for_for_asn_4568 , CONVOLUTION_LOOP_for_for_for_asn_4570});
  assign buf_acc_data_8_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4560
      , CONVOLUTION_LOOP_for_for_for_asn_4562 , CONVOLUTION_LOOP_for_for_for_asn_4564});
  assign buf_acc_data_8_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4554
      , CONVOLUTION_LOOP_for_for_for_asn_4556 , CONVOLUTION_LOOP_for_for_for_asn_4558});
  assign buf_acc_data_8_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4548
      , CONVOLUTION_LOOP_for_for_for_asn_4550 , CONVOLUTION_LOOP_for_for_for_asn_4552});
  assign buf_acc_data_8_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_8_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4542
      , CONVOLUTION_LOOP_for_for_for_asn_4544 , CONVOLUTION_LOOP_for_for_for_asn_4546});
  assign buf_acc_data_9_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4536
      , CONVOLUTION_LOOP_for_for_for_asn_4538 , CONVOLUTION_LOOP_for_for_for_asn_4540});
  assign buf_acc_data_9_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4530
      , CONVOLUTION_LOOP_for_for_for_asn_4532 , CONVOLUTION_LOOP_for_for_for_asn_4534});
  assign buf_acc_data_9_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4524
      , CONVOLUTION_LOOP_for_for_for_asn_4526 , CONVOLUTION_LOOP_for_for_for_asn_4528});
  assign buf_acc_data_9_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4518
      , CONVOLUTION_LOOP_for_for_for_asn_4520 , CONVOLUTION_LOOP_for_for_for_asn_4522});
  assign buf_acc_data_9_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4512
      , CONVOLUTION_LOOP_for_for_for_asn_4514 , CONVOLUTION_LOOP_for_for_for_asn_4516});
  assign buf_acc_data_9_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4506
      , CONVOLUTION_LOOP_for_for_for_asn_4508 , CONVOLUTION_LOOP_for_for_for_asn_4510});
  assign buf_acc_data_9_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4500
      , CONVOLUTION_LOOP_for_for_for_asn_4502 , CONVOLUTION_LOOP_for_for_for_asn_4504});
  assign buf_acc_data_9_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4494
      , CONVOLUTION_LOOP_for_for_for_asn_4496 , CONVOLUTION_LOOP_for_for_for_asn_4498});
  assign buf_acc_data_9_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4488
      , CONVOLUTION_LOOP_for_for_for_asn_4490 , CONVOLUTION_LOOP_for_for_for_asn_4492});
  assign buf_acc_data_9_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4482
      , CONVOLUTION_LOOP_for_for_for_asn_4484 , CONVOLUTION_LOOP_for_for_for_asn_4486});
  assign buf_acc_data_9_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4476
      , CONVOLUTION_LOOP_for_for_for_asn_4478 , CONVOLUTION_LOOP_for_for_for_asn_4480});
  assign buf_acc_data_9_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4470
      , CONVOLUTION_LOOP_for_for_for_asn_4472 , CONVOLUTION_LOOP_for_for_for_asn_4474});
  assign buf_acc_data_9_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4464
      , CONVOLUTION_LOOP_for_for_for_asn_4466 , CONVOLUTION_LOOP_for_for_for_asn_4468});
  assign buf_acc_data_9_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4458
      , CONVOLUTION_LOOP_for_for_for_asn_4460 , CONVOLUTION_LOOP_for_for_for_asn_4462});
  assign buf_acc_data_9_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4452
      , CONVOLUTION_LOOP_for_for_for_asn_4454 , CONVOLUTION_LOOP_for_for_for_asn_4456});
  assign buf_acc_data_9_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4446
      , CONVOLUTION_LOOP_for_for_for_asn_4448 , CONVOLUTION_LOOP_for_for_for_asn_4450});
  assign buf_acc_data_9_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4440
      , CONVOLUTION_LOOP_for_for_for_asn_4442 , CONVOLUTION_LOOP_for_for_for_asn_4444});
  assign buf_acc_data_9_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_9_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4434
      , CONVOLUTION_LOOP_for_for_for_asn_4436 , CONVOLUTION_LOOP_for_for_for_asn_4438});
  assign buf_acc_data_10_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4428
      , CONVOLUTION_LOOP_for_for_for_asn_4430 , CONVOLUTION_LOOP_for_for_for_asn_4432});
  assign buf_acc_data_10_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4422
      , CONVOLUTION_LOOP_for_for_for_asn_4424 , CONVOLUTION_LOOP_for_for_for_asn_4426});
  assign buf_acc_data_10_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4416
      , CONVOLUTION_LOOP_for_for_for_asn_4418 , CONVOLUTION_LOOP_for_for_for_asn_4420});
  assign buf_acc_data_10_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4410
      , CONVOLUTION_LOOP_for_for_for_asn_4412 , CONVOLUTION_LOOP_for_for_for_asn_4414});
  assign buf_acc_data_10_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4404
      , CONVOLUTION_LOOP_for_for_for_asn_4406 , CONVOLUTION_LOOP_for_for_for_asn_4408});
  assign buf_acc_data_10_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4398
      , CONVOLUTION_LOOP_for_for_for_asn_4400 , CONVOLUTION_LOOP_for_for_for_asn_4402});
  assign buf_acc_data_10_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4392
      , CONVOLUTION_LOOP_for_for_for_asn_4394 , CONVOLUTION_LOOP_for_for_for_asn_4396});
  assign buf_acc_data_10_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4386
      , CONVOLUTION_LOOP_for_for_for_asn_4388 , CONVOLUTION_LOOP_for_for_for_asn_4390});
  assign buf_acc_data_10_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4380
      , CONVOLUTION_LOOP_for_for_for_asn_4382 , CONVOLUTION_LOOP_for_for_for_asn_4384});
  assign buf_acc_data_10_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4374
      , CONVOLUTION_LOOP_for_for_for_asn_4376 , CONVOLUTION_LOOP_for_for_for_asn_4378});
  assign buf_acc_data_10_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4368
      , CONVOLUTION_LOOP_for_for_for_asn_4370 , CONVOLUTION_LOOP_for_for_for_asn_4372});
  assign buf_acc_data_10_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4362
      , CONVOLUTION_LOOP_for_for_for_asn_4364 , CONVOLUTION_LOOP_for_for_for_asn_4366});
  assign buf_acc_data_10_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4356
      , CONVOLUTION_LOOP_for_for_for_asn_4358 , CONVOLUTION_LOOP_for_for_for_asn_4360});
  assign buf_acc_data_10_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4350
      , CONVOLUTION_LOOP_for_for_for_asn_4352 , CONVOLUTION_LOOP_for_for_for_asn_4354});
  assign buf_acc_data_10_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4344
      , CONVOLUTION_LOOP_for_for_for_asn_4346 , CONVOLUTION_LOOP_for_for_for_asn_4348});
  assign buf_acc_data_10_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4338
      , CONVOLUTION_LOOP_for_for_for_asn_4340 , CONVOLUTION_LOOP_for_for_for_asn_4342});
  assign buf_acc_data_10_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4332
      , CONVOLUTION_LOOP_for_for_for_asn_4334 , CONVOLUTION_LOOP_for_for_for_asn_4336});
  assign buf_acc_data_10_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_10_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4326
      , CONVOLUTION_LOOP_for_for_for_asn_4328 , CONVOLUTION_LOOP_for_for_for_asn_4330});
  assign buf_acc_data_11_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4320
      , CONVOLUTION_LOOP_for_for_for_asn_4322 , CONVOLUTION_LOOP_for_for_for_asn_4324});
  assign buf_acc_data_11_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4314
      , CONVOLUTION_LOOP_for_for_for_asn_4316 , CONVOLUTION_LOOP_for_for_for_asn_4318});
  assign buf_acc_data_11_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4308
      , CONVOLUTION_LOOP_for_for_for_asn_4310 , CONVOLUTION_LOOP_for_for_for_asn_4312});
  assign buf_acc_data_11_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4302
      , CONVOLUTION_LOOP_for_for_for_asn_4304 , CONVOLUTION_LOOP_for_for_for_asn_4306});
  assign buf_acc_data_11_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4296
      , CONVOLUTION_LOOP_for_for_for_asn_4298 , CONVOLUTION_LOOP_for_for_for_asn_4300});
  assign buf_acc_data_11_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4290
      , CONVOLUTION_LOOP_for_for_for_asn_4292 , CONVOLUTION_LOOP_for_for_for_asn_4294});
  assign buf_acc_data_11_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4284
      , CONVOLUTION_LOOP_for_for_for_asn_4286 , CONVOLUTION_LOOP_for_for_for_asn_4288});
  assign buf_acc_data_11_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4278
      , CONVOLUTION_LOOP_for_for_for_asn_4280 , CONVOLUTION_LOOP_for_for_for_asn_4282});
  assign buf_acc_data_11_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4272
      , CONVOLUTION_LOOP_for_for_for_asn_4274 , CONVOLUTION_LOOP_for_for_for_asn_4276});
  assign buf_acc_data_11_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4266
      , CONVOLUTION_LOOP_for_for_for_asn_4268 , CONVOLUTION_LOOP_for_for_for_asn_4270});
  assign buf_acc_data_11_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4260
      , CONVOLUTION_LOOP_for_for_for_asn_4262 , CONVOLUTION_LOOP_for_for_for_asn_4264});
  assign buf_acc_data_11_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4254
      , CONVOLUTION_LOOP_for_for_for_asn_4256 , CONVOLUTION_LOOP_for_for_for_asn_4258});
  assign buf_acc_data_11_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4248
      , CONVOLUTION_LOOP_for_for_for_asn_4250 , CONVOLUTION_LOOP_for_for_for_asn_4252});
  assign buf_acc_data_11_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4242
      , CONVOLUTION_LOOP_for_for_for_asn_4244 , CONVOLUTION_LOOP_for_for_for_asn_4246});
  assign buf_acc_data_11_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4236
      , CONVOLUTION_LOOP_for_for_for_asn_4238 , CONVOLUTION_LOOP_for_for_for_asn_4240});
  assign buf_acc_data_11_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4230
      , CONVOLUTION_LOOP_for_for_for_asn_4232 , CONVOLUTION_LOOP_for_for_for_asn_4234});
  assign buf_acc_data_11_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4224
      , CONVOLUTION_LOOP_for_for_for_asn_4226 , CONVOLUTION_LOOP_for_for_for_asn_4228});
  assign buf_acc_data_11_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_11_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4218
      , CONVOLUTION_LOOP_for_for_for_asn_4220 , CONVOLUTION_LOOP_for_for_for_asn_4222});
  assign buf_acc_data_12_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4212
      , CONVOLUTION_LOOP_for_for_for_asn_4214 , CONVOLUTION_LOOP_for_for_for_asn_4216});
  assign buf_acc_data_12_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4206
      , CONVOLUTION_LOOP_for_for_for_asn_4208 , CONVOLUTION_LOOP_for_for_for_asn_4210});
  assign buf_acc_data_12_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4200
      , CONVOLUTION_LOOP_for_for_for_asn_4202 , CONVOLUTION_LOOP_for_for_for_asn_4204});
  assign buf_acc_data_12_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4194
      , CONVOLUTION_LOOP_for_for_for_asn_4196 , CONVOLUTION_LOOP_for_for_for_asn_4198});
  assign buf_acc_data_12_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4188
      , CONVOLUTION_LOOP_for_for_for_asn_4190 , CONVOLUTION_LOOP_for_for_for_asn_4192});
  assign buf_acc_data_12_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4182
      , CONVOLUTION_LOOP_for_for_for_asn_4184 , CONVOLUTION_LOOP_for_for_for_asn_4186});
  assign buf_acc_data_12_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4176
      , CONVOLUTION_LOOP_for_for_for_asn_4178 , CONVOLUTION_LOOP_for_for_for_asn_4180});
  assign buf_acc_data_12_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4170
      , CONVOLUTION_LOOP_for_for_for_asn_4172 , CONVOLUTION_LOOP_for_for_for_asn_4174});
  assign buf_acc_data_12_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4164
      , CONVOLUTION_LOOP_for_for_for_asn_4166 , CONVOLUTION_LOOP_for_for_for_asn_4168});
  assign buf_acc_data_12_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4158
      , CONVOLUTION_LOOP_for_for_for_asn_4160 , CONVOLUTION_LOOP_for_for_for_asn_4162});
  assign buf_acc_data_12_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4152
      , CONVOLUTION_LOOP_for_for_for_asn_4154 , CONVOLUTION_LOOP_for_for_for_asn_4156});
  assign buf_acc_data_12_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4146
      , CONVOLUTION_LOOP_for_for_for_asn_4148 , CONVOLUTION_LOOP_for_for_for_asn_4150});
  assign buf_acc_data_12_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4140
      , CONVOLUTION_LOOP_for_for_for_asn_4142 , CONVOLUTION_LOOP_for_for_for_asn_4144});
  assign buf_acc_data_12_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4134
      , CONVOLUTION_LOOP_for_for_for_asn_4136 , CONVOLUTION_LOOP_for_for_for_asn_4138});
  assign buf_acc_data_12_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4128
      , CONVOLUTION_LOOP_for_for_for_asn_4130 , CONVOLUTION_LOOP_for_for_for_asn_4132});
  assign buf_acc_data_12_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4122
      , CONVOLUTION_LOOP_for_for_for_asn_4124 , CONVOLUTION_LOOP_for_for_for_asn_4126});
  assign buf_acc_data_12_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4116
      , CONVOLUTION_LOOP_for_for_for_asn_4118 , CONVOLUTION_LOOP_for_for_for_asn_4120});
  assign buf_acc_data_12_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_12_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4110
      , CONVOLUTION_LOOP_for_for_for_asn_4112 , CONVOLUTION_LOOP_for_for_for_asn_4114});
  assign buf_acc_data_13_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4104
      , CONVOLUTION_LOOP_for_for_for_asn_4106 , CONVOLUTION_LOOP_for_for_for_asn_4108});
  assign buf_acc_data_13_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4098
      , CONVOLUTION_LOOP_for_for_for_asn_4100 , CONVOLUTION_LOOP_for_for_for_asn_4102});
  assign buf_acc_data_13_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4092
      , CONVOLUTION_LOOP_for_for_for_asn_4094 , CONVOLUTION_LOOP_for_for_for_asn_4096});
  assign buf_acc_data_13_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4086
      , CONVOLUTION_LOOP_for_for_for_asn_4088 , CONVOLUTION_LOOP_for_for_for_asn_4090});
  assign buf_acc_data_13_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4080
      , CONVOLUTION_LOOP_for_for_for_asn_4082 , CONVOLUTION_LOOP_for_for_for_asn_4084});
  assign buf_acc_data_13_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4074
      , CONVOLUTION_LOOP_for_for_for_asn_4076 , CONVOLUTION_LOOP_for_for_for_asn_4078});
  assign buf_acc_data_13_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4068
      , CONVOLUTION_LOOP_for_for_for_asn_4070 , CONVOLUTION_LOOP_for_for_for_asn_4072});
  assign buf_acc_data_13_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4062
      , CONVOLUTION_LOOP_for_for_for_asn_4064 , CONVOLUTION_LOOP_for_for_for_asn_4066});
  assign buf_acc_data_13_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4056
      , CONVOLUTION_LOOP_for_for_for_asn_4058 , CONVOLUTION_LOOP_for_for_for_asn_4060});
  assign buf_acc_data_13_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4050
      , CONVOLUTION_LOOP_for_for_for_asn_4052 , CONVOLUTION_LOOP_for_for_for_asn_4054});
  assign buf_acc_data_13_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4044
      , CONVOLUTION_LOOP_for_for_for_asn_4046 , CONVOLUTION_LOOP_for_for_for_asn_4048});
  assign buf_acc_data_13_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4038
      , CONVOLUTION_LOOP_for_for_for_asn_4040 , CONVOLUTION_LOOP_for_for_for_asn_4042});
  assign buf_acc_data_13_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4032
      , CONVOLUTION_LOOP_for_for_for_asn_4034 , CONVOLUTION_LOOP_for_for_for_asn_4036});
  assign buf_acc_data_13_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4026
      , CONVOLUTION_LOOP_for_for_for_asn_4028 , CONVOLUTION_LOOP_for_for_for_asn_4030});
  assign buf_acc_data_13_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4020
      , CONVOLUTION_LOOP_for_for_for_asn_4022 , CONVOLUTION_LOOP_for_for_for_asn_4024});
  assign buf_acc_data_13_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4014
      , CONVOLUTION_LOOP_for_for_for_asn_4016 , CONVOLUTION_LOOP_for_for_for_asn_4018});
  assign buf_acc_data_13_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4008
      , CONVOLUTION_LOOP_for_for_for_asn_4010 , CONVOLUTION_LOOP_for_for_for_asn_4012});
  assign buf_acc_data_13_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_13_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4002
      , CONVOLUTION_LOOP_for_for_for_asn_4004 , CONVOLUTION_LOOP_for_for_for_asn_4006});
  assign buf_acc_data_14_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3996
      , CONVOLUTION_LOOP_for_for_for_asn_3998 , CONVOLUTION_LOOP_for_for_for_asn_4000});
  assign buf_acc_data_14_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3990
      , CONVOLUTION_LOOP_for_for_for_asn_3992 , CONVOLUTION_LOOP_for_for_for_asn_3994});
  assign buf_acc_data_14_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3984
      , CONVOLUTION_LOOP_for_for_for_asn_3986 , CONVOLUTION_LOOP_for_for_for_asn_3988});
  assign buf_acc_data_14_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3978
      , CONVOLUTION_LOOP_for_for_for_asn_3980 , CONVOLUTION_LOOP_for_for_for_asn_3982});
  assign buf_acc_data_14_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3972
      , CONVOLUTION_LOOP_for_for_for_asn_3974 , CONVOLUTION_LOOP_for_for_for_asn_3976});
  assign buf_acc_data_14_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3966
      , CONVOLUTION_LOOP_for_for_for_asn_3968 , CONVOLUTION_LOOP_for_for_for_asn_3970});
  assign buf_acc_data_14_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3960
      , CONVOLUTION_LOOP_for_for_for_asn_3962 , CONVOLUTION_LOOP_for_for_for_asn_3964});
  assign buf_acc_data_14_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3954
      , CONVOLUTION_LOOP_for_for_for_asn_3956 , CONVOLUTION_LOOP_for_for_for_asn_3958});
  assign buf_acc_data_14_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3948
      , CONVOLUTION_LOOP_for_for_for_asn_3950 , CONVOLUTION_LOOP_for_for_for_asn_3952});
  assign buf_acc_data_14_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3942
      , CONVOLUTION_LOOP_for_for_for_asn_3944 , CONVOLUTION_LOOP_for_for_for_asn_3946});
  assign buf_acc_data_14_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3936
      , CONVOLUTION_LOOP_for_for_for_asn_3938 , CONVOLUTION_LOOP_for_for_for_asn_3940});
  assign buf_acc_data_14_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3930
      , CONVOLUTION_LOOP_for_for_for_asn_3932 , CONVOLUTION_LOOP_for_for_for_asn_3934});
  assign buf_acc_data_14_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3924
      , CONVOLUTION_LOOP_for_for_for_asn_3926 , CONVOLUTION_LOOP_for_for_for_asn_3928});
  assign buf_acc_data_14_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3918
      , CONVOLUTION_LOOP_for_for_for_asn_3920 , CONVOLUTION_LOOP_for_for_for_asn_3922});
  assign buf_acc_data_14_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3912
      , CONVOLUTION_LOOP_for_for_for_asn_3914 , CONVOLUTION_LOOP_for_for_for_asn_3916});
  assign buf_acc_data_14_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3906
      , CONVOLUTION_LOOP_for_for_for_asn_3908 , CONVOLUTION_LOOP_for_for_for_asn_3910});
  assign buf_acc_data_14_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3900
      , CONVOLUTION_LOOP_for_for_for_asn_3902 , CONVOLUTION_LOOP_for_for_for_asn_3904});
  assign buf_acc_data_14_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_14_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3894
      , CONVOLUTION_LOOP_for_for_for_asn_3896 , CONVOLUTION_LOOP_for_for_for_asn_3898});
  assign buf_acc_data_15_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3888
      , CONVOLUTION_LOOP_for_for_for_asn_3890 , CONVOLUTION_LOOP_for_for_for_asn_3892});
  assign buf_acc_data_15_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3882
      , CONVOLUTION_LOOP_for_for_for_asn_3884 , CONVOLUTION_LOOP_for_for_for_asn_3886});
  assign buf_acc_data_15_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3876
      , CONVOLUTION_LOOP_for_for_for_asn_3878 , CONVOLUTION_LOOP_for_for_for_asn_3880});
  assign buf_acc_data_15_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3870
      , CONVOLUTION_LOOP_for_for_for_asn_3872 , CONVOLUTION_LOOP_for_for_for_asn_3874});
  assign buf_acc_data_15_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3864
      , CONVOLUTION_LOOP_for_for_for_asn_3866 , CONVOLUTION_LOOP_for_for_for_asn_3868});
  assign buf_acc_data_15_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3858
      , CONVOLUTION_LOOP_for_for_for_asn_3860 , CONVOLUTION_LOOP_for_for_for_asn_3862});
  assign buf_acc_data_15_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3852
      , CONVOLUTION_LOOP_for_for_for_asn_3854 , CONVOLUTION_LOOP_for_for_for_asn_3856});
  assign buf_acc_data_15_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3846
      , CONVOLUTION_LOOP_for_for_for_asn_3848 , CONVOLUTION_LOOP_for_for_for_asn_3850});
  assign buf_acc_data_15_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3840
      , CONVOLUTION_LOOP_for_for_for_asn_3842 , CONVOLUTION_LOOP_for_for_for_asn_3844});
  assign buf_acc_data_15_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3834
      , CONVOLUTION_LOOP_for_for_for_asn_3836 , CONVOLUTION_LOOP_for_for_for_asn_3838});
  assign buf_acc_data_15_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3828
      , CONVOLUTION_LOOP_for_for_for_asn_3830 , CONVOLUTION_LOOP_for_for_for_asn_3832});
  assign buf_acc_data_15_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3822
      , CONVOLUTION_LOOP_for_for_for_asn_3824 , CONVOLUTION_LOOP_for_for_for_asn_3826});
  assign buf_acc_data_15_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3816
      , CONVOLUTION_LOOP_for_for_for_asn_3818 , CONVOLUTION_LOOP_for_for_for_asn_3820});
  assign buf_acc_data_15_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3810
      , CONVOLUTION_LOOP_for_for_for_asn_3812 , CONVOLUTION_LOOP_for_for_for_asn_3814});
  assign buf_acc_data_15_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3804
      , CONVOLUTION_LOOP_for_for_for_asn_3806 , CONVOLUTION_LOOP_for_for_for_asn_3808});
  assign buf_acc_data_15_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3798
      , CONVOLUTION_LOOP_for_for_for_asn_3800 , CONVOLUTION_LOOP_for_for_for_asn_3802});
  assign buf_acc_data_15_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3792
      , CONVOLUTION_LOOP_for_for_for_asn_3794 , CONVOLUTION_LOOP_for_for_for_asn_3796});
  assign buf_acc_data_15_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_15_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3786
      , CONVOLUTION_LOOP_for_for_for_asn_3788 , CONVOLUTION_LOOP_for_for_for_asn_3790});
  assign buf_acc_data_16_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3780
      , CONVOLUTION_LOOP_for_for_for_asn_3782 , CONVOLUTION_LOOP_for_for_for_asn_3784});
  assign buf_acc_data_16_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3774
      , CONVOLUTION_LOOP_for_for_for_asn_3776 , CONVOLUTION_LOOP_for_for_for_asn_3778});
  assign buf_acc_data_16_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3768
      , CONVOLUTION_LOOP_for_for_for_asn_3770 , CONVOLUTION_LOOP_for_for_for_asn_3772});
  assign buf_acc_data_16_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3762
      , CONVOLUTION_LOOP_for_for_for_asn_3764 , CONVOLUTION_LOOP_for_for_for_asn_3766});
  assign buf_acc_data_16_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3756
      , CONVOLUTION_LOOP_for_for_for_asn_3758 , CONVOLUTION_LOOP_for_for_for_asn_3760});
  assign buf_acc_data_16_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3750
      , CONVOLUTION_LOOP_for_for_for_asn_3752 , CONVOLUTION_LOOP_for_for_for_asn_3754});
  assign buf_acc_data_16_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3744
      , CONVOLUTION_LOOP_for_for_for_asn_3746 , CONVOLUTION_LOOP_for_for_for_asn_3748});
  assign buf_acc_data_16_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3738
      , CONVOLUTION_LOOP_for_for_for_asn_3740 , CONVOLUTION_LOOP_for_for_for_asn_3742});
  assign buf_acc_data_16_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3732
      , CONVOLUTION_LOOP_for_for_for_asn_3734 , CONVOLUTION_LOOP_for_for_for_asn_3736});
  assign buf_acc_data_16_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3726
      , CONVOLUTION_LOOP_for_for_for_asn_3728 , CONVOLUTION_LOOP_for_for_for_asn_3730});
  assign buf_acc_data_16_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3720
      , CONVOLUTION_LOOP_for_for_for_asn_3722 , CONVOLUTION_LOOP_for_for_for_asn_3724});
  assign buf_acc_data_16_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3714
      , CONVOLUTION_LOOP_for_for_for_asn_3716 , CONVOLUTION_LOOP_for_for_for_asn_3718});
  assign buf_acc_data_16_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3708
      , CONVOLUTION_LOOP_for_for_for_asn_3710 , CONVOLUTION_LOOP_for_for_for_asn_3712});
  assign buf_acc_data_16_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3702
      , CONVOLUTION_LOOP_for_for_for_asn_3704 , CONVOLUTION_LOOP_for_for_for_asn_3706});
  assign buf_acc_data_16_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3696
      , CONVOLUTION_LOOP_for_for_for_asn_3698 , CONVOLUTION_LOOP_for_for_for_asn_3700});
  assign buf_acc_data_16_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3690
      , CONVOLUTION_LOOP_for_for_for_asn_3692 , CONVOLUTION_LOOP_for_for_for_asn_3694});
  assign buf_acc_data_16_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3684
      , CONVOLUTION_LOOP_for_for_for_asn_3686 , CONVOLUTION_LOOP_for_for_for_asn_3688});
  assign buf_acc_data_16_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_16_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3678
      , CONVOLUTION_LOOP_for_for_for_asn_3680 , CONVOLUTION_LOOP_for_for_for_asn_3682});
  assign buf_acc_data_17_0_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_0_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3672
      , CONVOLUTION_LOOP_for_for_for_asn_3674 , CONVOLUTION_LOOP_for_for_for_asn_3676});
  assign buf_acc_data_17_1_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_1_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3666
      , CONVOLUTION_LOOP_for_for_for_asn_3668 , CONVOLUTION_LOOP_for_for_for_asn_3670});
  assign buf_acc_data_17_2_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_2_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3660
      , CONVOLUTION_LOOP_for_for_for_asn_3662 , CONVOLUTION_LOOP_for_for_for_asn_3664});
  assign buf_acc_data_17_3_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_3_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3654
      , CONVOLUTION_LOOP_for_for_for_asn_3656 , CONVOLUTION_LOOP_for_for_for_asn_3658});
  assign buf_acc_data_17_4_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_4_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3648
      , CONVOLUTION_LOOP_for_for_for_asn_3650 , CONVOLUTION_LOOP_for_for_for_asn_3652});
  assign buf_acc_data_17_5_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_5_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3642
      , CONVOLUTION_LOOP_for_for_for_asn_3644 , CONVOLUTION_LOOP_for_for_for_asn_3646});
  assign buf_acc_data_17_6_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_6_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3636
      , CONVOLUTION_LOOP_for_for_for_asn_3638 , CONVOLUTION_LOOP_for_for_for_asn_3640});
  assign buf_acc_data_17_7_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_7_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3630
      , CONVOLUTION_LOOP_for_for_for_asn_3632 , CONVOLUTION_LOOP_for_for_for_asn_3634});
  assign buf_acc_data_17_8_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_8_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3624
      , CONVOLUTION_LOOP_for_for_for_asn_3626 , CONVOLUTION_LOOP_for_for_for_asn_3628});
  assign buf_acc_data_17_9_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_9_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3618
      , CONVOLUTION_LOOP_for_for_for_asn_3620 , CONVOLUTION_LOOP_for_for_for_asn_3622});
  assign buf_acc_data_17_10_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_10_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3612
      , CONVOLUTION_LOOP_for_for_for_asn_3614 , CONVOLUTION_LOOP_for_for_for_asn_3616});
  assign buf_acc_data_17_11_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_11_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3606
      , CONVOLUTION_LOOP_for_for_for_asn_3608 , CONVOLUTION_LOOP_for_for_for_asn_3610});
  assign buf_acc_data_17_12_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_12_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3600
      , CONVOLUTION_LOOP_for_for_for_asn_3602 , CONVOLUTION_LOOP_for_for_for_asn_3604});
  assign buf_acc_data_17_13_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_13_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3594
      , CONVOLUTION_LOOP_for_for_for_asn_3596 , CONVOLUTION_LOOP_for_for_for_asn_3598});
  assign buf_acc_data_17_14_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_14_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3588
      , CONVOLUTION_LOOP_for_for_for_asn_3590 , CONVOLUTION_LOOP_for_for_for_asn_3592});
  assign buf_acc_data_17_15_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_15_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3582
      , CONVOLUTION_LOOP_for_for_for_asn_3584 , CONVOLUTION_LOOP_for_for_for_asn_3586});
  assign buf_acc_data_17_16_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_16_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3576
      , CONVOLUTION_LOOP_for_for_for_asn_3578 , CONVOLUTION_LOOP_for_for_for_asn_3580});
  assign buf_acc_data_17_17_56_46_sva_dfm_1 = MUX1HOT_v_11_3_2(buf_acc_data_17_17_56_46_sva,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_2}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3570
      , CONVOLUTION_LOOP_for_for_for_asn_3572 , CONVOLUTION_LOOP_for_for_for_asn_3574});
  assign buf_acc_data_0_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5508 , CONVOLUTION_LOOP_for_for_for_asn_5510
      , CONVOLUTION_LOOP_for_for_for_asn_5512});
  assign buf_acc_data_0_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5502 , CONVOLUTION_LOOP_for_for_for_asn_5504
      , CONVOLUTION_LOOP_for_for_for_asn_5506});
  assign buf_acc_data_0_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5496 , CONVOLUTION_LOOP_for_for_for_asn_5498
      , CONVOLUTION_LOOP_for_for_for_asn_5500});
  assign buf_acc_data_0_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5490 , CONVOLUTION_LOOP_for_for_for_asn_5492
      , CONVOLUTION_LOOP_for_for_for_asn_5494});
  assign buf_acc_data_0_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5484 , CONVOLUTION_LOOP_for_for_for_asn_5486
      , CONVOLUTION_LOOP_for_for_for_asn_5488});
  assign buf_acc_data_0_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5478 , CONVOLUTION_LOOP_for_for_for_asn_5480
      , CONVOLUTION_LOOP_for_for_for_asn_5482});
  assign buf_acc_data_0_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5472 , CONVOLUTION_LOOP_for_for_for_asn_5474
      , CONVOLUTION_LOOP_for_for_for_asn_5476});
  assign buf_acc_data_0_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5466 , CONVOLUTION_LOOP_for_for_for_asn_5468
      , CONVOLUTION_LOOP_for_for_for_asn_5470});
  assign buf_acc_data_0_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5460 , CONVOLUTION_LOOP_for_for_for_asn_5462
      , CONVOLUTION_LOOP_for_for_for_asn_5464});
  assign buf_acc_data_0_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5454 , CONVOLUTION_LOOP_for_for_for_asn_5456
      , CONVOLUTION_LOOP_for_for_for_asn_5458});
  assign buf_acc_data_0_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5448 , CONVOLUTION_LOOP_for_for_for_asn_5450
      , CONVOLUTION_LOOP_for_for_for_asn_5452});
  assign buf_acc_data_0_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5442 , CONVOLUTION_LOOP_for_for_for_asn_5444
      , CONVOLUTION_LOOP_for_for_for_asn_5446});
  assign buf_acc_data_0_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5436 , CONVOLUTION_LOOP_for_for_for_asn_5438
      , CONVOLUTION_LOOP_for_for_for_asn_5440});
  assign buf_acc_data_0_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5430 , CONVOLUTION_LOOP_for_for_for_asn_5432
      , CONVOLUTION_LOOP_for_for_for_asn_5434});
  assign buf_acc_data_0_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5424 , CONVOLUTION_LOOP_for_for_for_asn_5426
      , CONVOLUTION_LOOP_for_for_for_asn_5428});
  assign buf_acc_data_0_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5418 , CONVOLUTION_LOOP_for_for_for_asn_5420
      , CONVOLUTION_LOOP_for_for_for_asn_5422});
  assign buf_acc_data_0_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5412 , CONVOLUTION_LOOP_for_for_for_asn_5414
      , CONVOLUTION_LOOP_for_for_for_asn_5416});
  assign buf_acc_data_0_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_0_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5406 , CONVOLUTION_LOOP_for_for_for_asn_5408
      , CONVOLUTION_LOOP_for_for_for_asn_5410});
  assign buf_acc_data_1_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5400 , CONVOLUTION_LOOP_for_for_for_asn_5402
      , CONVOLUTION_LOOP_for_for_for_asn_5404});
  assign buf_acc_data_1_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5394 , CONVOLUTION_LOOP_for_for_for_asn_5396
      , CONVOLUTION_LOOP_for_for_for_asn_5398});
  assign buf_acc_data_1_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5388 , CONVOLUTION_LOOP_for_for_for_asn_5390
      , CONVOLUTION_LOOP_for_for_for_asn_5392});
  assign buf_acc_data_1_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5382 , CONVOLUTION_LOOP_for_for_for_asn_5384
      , CONVOLUTION_LOOP_for_for_for_asn_5386});
  assign buf_acc_data_1_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5376 , CONVOLUTION_LOOP_for_for_for_asn_5378
      , CONVOLUTION_LOOP_for_for_for_asn_5380});
  assign buf_acc_data_1_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5370 , CONVOLUTION_LOOP_for_for_for_asn_5372
      , CONVOLUTION_LOOP_for_for_for_asn_5374});
  assign buf_acc_data_1_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5364 , CONVOLUTION_LOOP_for_for_for_asn_5366
      , CONVOLUTION_LOOP_for_for_for_asn_5368});
  assign buf_acc_data_1_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5358 , CONVOLUTION_LOOP_for_for_for_asn_5360
      , CONVOLUTION_LOOP_for_for_for_asn_5362});
  assign buf_acc_data_1_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5352 , CONVOLUTION_LOOP_for_for_for_asn_5354
      , CONVOLUTION_LOOP_for_for_for_asn_5356});
  assign buf_acc_data_1_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5346 , CONVOLUTION_LOOP_for_for_for_asn_5348
      , CONVOLUTION_LOOP_for_for_for_asn_5350});
  assign buf_acc_data_1_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5340 , CONVOLUTION_LOOP_for_for_for_asn_5342
      , CONVOLUTION_LOOP_for_for_for_asn_5344});
  assign buf_acc_data_1_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5334 , CONVOLUTION_LOOP_for_for_for_asn_5336
      , CONVOLUTION_LOOP_for_for_for_asn_5338});
  assign buf_acc_data_1_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5328 , CONVOLUTION_LOOP_for_for_for_asn_5330
      , CONVOLUTION_LOOP_for_for_for_asn_5332});
  assign buf_acc_data_1_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5322 , CONVOLUTION_LOOP_for_for_for_asn_5324
      , CONVOLUTION_LOOP_for_for_for_asn_5326});
  assign buf_acc_data_1_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5316 , CONVOLUTION_LOOP_for_for_for_asn_5318
      , CONVOLUTION_LOOP_for_for_for_asn_5320});
  assign buf_acc_data_1_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5310 , CONVOLUTION_LOOP_for_for_for_asn_5312
      , CONVOLUTION_LOOP_for_for_for_asn_5314});
  assign buf_acc_data_1_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5304 , CONVOLUTION_LOOP_for_for_for_asn_5306
      , CONVOLUTION_LOOP_for_for_for_asn_5308});
  assign buf_acc_data_1_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_1_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5298 , CONVOLUTION_LOOP_for_for_for_asn_5300
      , CONVOLUTION_LOOP_for_for_for_asn_5302});
  assign buf_acc_data_2_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5292 , CONVOLUTION_LOOP_for_for_for_asn_5294
      , CONVOLUTION_LOOP_for_for_for_asn_5296});
  assign buf_acc_data_2_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5286 , CONVOLUTION_LOOP_for_for_for_asn_5288
      , CONVOLUTION_LOOP_for_for_for_asn_5290});
  assign buf_acc_data_2_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5280 , CONVOLUTION_LOOP_for_for_for_asn_5282
      , CONVOLUTION_LOOP_for_for_for_asn_5284});
  assign buf_acc_data_2_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5274 , CONVOLUTION_LOOP_for_for_for_asn_5276
      , CONVOLUTION_LOOP_for_for_for_asn_5278});
  assign buf_acc_data_2_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5268 , CONVOLUTION_LOOP_for_for_for_asn_5270
      , CONVOLUTION_LOOP_for_for_for_asn_5272});
  assign buf_acc_data_2_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5262 , CONVOLUTION_LOOP_for_for_for_asn_5264
      , CONVOLUTION_LOOP_for_for_for_asn_5266});
  assign buf_acc_data_2_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5256 , CONVOLUTION_LOOP_for_for_for_asn_5258
      , CONVOLUTION_LOOP_for_for_for_asn_5260});
  assign buf_acc_data_2_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5250 , CONVOLUTION_LOOP_for_for_for_asn_5252
      , CONVOLUTION_LOOP_for_for_for_asn_5254});
  assign buf_acc_data_2_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5244 , CONVOLUTION_LOOP_for_for_for_asn_5246
      , CONVOLUTION_LOOP_for_for_for_asn_5248});
  assign buf_acc_data_2_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5238 , CONVOLUTION_LOOP_for_for_for_asn_5240
      , CONVOLUTION_LOOP_for_for_for_asn_5242});
  assign buf_acc_data_2_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5232 , CONVOLUTION_LOOP_for_for_for_asn_5234
      , CONVOLUTION_LOOP_for_for_for_asn_5236});
  assign buf_acc_data_2_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5226 , CONVOLUTION_LOOP_for_for_for_asn_5228
      , CONVOLUTION_LOOP_for_for_for_asn_5230});
  assign buf_acc_data_2_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5220 , CONVOLUTION_LOOP_for_for_for_asn_5222
      , CONVOLUTION_LOOP_for_for_for_asn_5224});
  assign buf_acc_data_2_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5214 , CONVOLUTION_LOOP_for_for_for_asn_5216
      , CONVOLUTION_LOOP_for_for_for_asn_5218});
  assign buf_acc_data_2_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5208 , CONVOLUTION_LOOP_for_for_for_asn_5210
      , CONVOLUTION_LOOP_for_for_for_asn_5212});
  assign buf_acc_data_2_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5202 , CONVOLUTION_LOOP_for_for_for_asn_5204
      , CONVOLUTION_LOOP_for_for_for_asn_5206});
  assign buf_acc_data_2_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5196 , CONVOLUTION_LOOP_for_for_for_asn_5198
      , CONVOLUTION_LOOP_for_for_for_asn_5200});
  assign buf_acc_data_2_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_2_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5190 , CONVOLUTION_LOOP_for_for_for_asn_5192
      , CONVOLUTION_LOOP_for_for_for_asn_5194});
  assign buf_acc_data_3_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5184 , CONVOLUTION_LOOP_for_for_for_asn_5186
      , CONVOLUTION_LOOP_for_for_for_asn_5188});
  assign buf_acc_data_3_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5178 , CONVOLUTION_LOOP_for_for_for_asn_5180
      , CONVOLUTION_LOOP_for_for_for_asn_5182});
  assign buf_acc_data_3_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5172 , CONVOLUTION_LOOP_for_for_for_asn_5174
      , CONVOLUTION_LOOP_for_for_for_asn_5176});
  assign buf_acc_data_3_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5166 , CONVOLUTION_LOOP_for_for_for_asn_5168
      , CONVOLUTION_LOOP_for_for_for_asn_5170});
  assign buf_acc_data_3_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5160 , CONVOLUTION_LOOP_for_for_for_asn_5162
      , CONVOLUTION_LOOP_for_for_for_asn_5164});
  assign buf_acc_data_3_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5154 , CONVOLUTION_LOOP_for_for_for_asn_5156
      , CONVOLUTION_LOOP_for_for_for_asn_5158});
  assign buf_acc_data_3_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5148 , CONVOLUTION_LOOP_for_for_for_asn_5150
      , CONVOLUTION_LOOP_for_for_for_asn_5152});
  assign buf_acc_data_3_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5142 , CONVOLUTION_LOOP_for_for_for_asn_5144
      , CONVOLUTION_LOOP_for_for_for_asn_5146});
  assign buf_acc_data_3_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5136 , CONVOLUTION_LOOP_for_for_for_asn_5138
      , CONVOLUTION_LOOP_for_for_for_asn_5140});
  assign buf_acc_data_3_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5130 , CONVOLUTION_LOOP_for_for_for_asn_5132
      , CONVOLUTION_LOOP_for_for_for_asn_5134});
  assign buf_acc_data_3_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5124 , CONVOLUTION_LOOP_for_for_for_asn_5126
      , CONVOLUTION_LOOP_for_for_for_asn_5128});
  assign buf_acc_data_3_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5118 , CONVOLUTION_LOOP_for_for_for_asn_5120
      , CONVOLUTION_LOOP_for_for_for_asn_5122});
  assign buf_acc_data_3_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5112 , CONVOLUTION_LOOP_for_for_for_asn_5114
      , CONVOLUTION_LOOP_for_for_for_asn_5116});
  assign buf_acc_data_3_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5106 , CONVOLUTION_LOOP_for_for_for_asn_5108
      , CONVOLUTION_LOOP_for_for_for_asn_5110});
  assign buf_acc_data_3_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5100 , CONVOLUTION_LOOP_for_for_for_asn_5102
      , CONVOLUTION_LOOP_for_for_for_asn_5104});
  assign buf_acc_data_3_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5094 , CONVOLUTION_LOOP_for_for_for_asn_5096
      , CONVOLUTION_LOOP_for_for_for_asn_5098});
  assign buf_acc_data_3_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5088 , CONVOLUTION_LOOP_for_for_for_asn_5090
      , CONVOLUTION_LOOP_for_for_for_asn_5092});
  assign buf_acc_data_3_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_3_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5082 , CONVOLUTION_LOOP_for_for_for_asn_5084
      , CONVOLUTION_LOOP_for_for_for_asn_5086});
  assign buf_acc_data_4_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5076 , CONVOLUTION_LOOP_for_for_for_asn_5078
      , CONVOLUTION_LOOP_for_for_for_asn_5080});
  assign buf_acc_data_4_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5070 , CONVOLUTION_LOOP_for_for_for_asn_5072
      , CONVOLUTION_LOOP_for_for_for_asn_5074});
  assign buf_acc_data_4_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5064 , CONVOLUTION_LOOP_for_for_for_asn_5066
      , CONVOLUTION_LOOP_for_for_for_asn_5068});
  assign buf_acc_data_4_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5058 , CONVOLUTION_LOOP_for_for_for_asn_5060
      , CONVOLUTION_LOOP_for_for_for_asn_5062});
  assign buf_acc_data_4_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5052 , CONVOLUTION_LOOP_for_for_for_asn_5054
      , CONVOLUTION_LOOP_for_for_for_asn_5056});
  assign buf_acc_data_4_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5046 , CONVOLUTION_LOOP_for_for_for_asn_5048
      , CONVOLUTION_LOOP_for_for_for_asn_5050});
  assign buf_acc_data_4_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5040 , CONVOLUTION_LOOP_for_for_for_asn_5042
      , CONVOLUTION_LOOP_for_for_for_asn_5044});
  assign buf_acc_data_4_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5034 , CONVOLUTION_LOOP_for_for_for_asn_5036
      , CONVOLUTION_LOOP_for_for_for_asn_5038});
  assign buf_acc_data_4_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5028 , CONVOLUTION_LOOP_for_for_for_asn_5030
      , CONVOLUTION_LOOP_for_for_for_asn_5032});
  assign buf_acc_data_4_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5022 , CONVOLUTION_LOOP_for_for_for_asn_5024
      , CONVOLUTION_LOOP_for_for_for_asn_5026});
  assign buf_acc_data_4_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5016 , CONVOLUTION_LOOP_for_for_for_asn_5018
      , CONVOLUTION_LOOP_for_for_for_asn_5020});
  assign buf_acc_data_4_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5010 , CONVOLUTION_LOOP_for_for_for_asn_5012
      , CONVOLUTION_LOOP_for_for_for_asn_5014});
  assign buf_acc_data_4_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5004 , CONVOLUTION_LOOP_for_for_for_asn_5006
      , CONVOLUTION_LOOP_for_for_for_asn_5008});
  assign buf_acc_data_4_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4998 , CONVOLUTION_LOOP_for_for_for_asn_5000
      , CONVOLUTION_LOOP_for_for_for_asn_5002});
  assign buf_acc_data_4_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4992 , CONVOLUTION_LOOP_for_for_for_asn_4994
      , CONVOLUTION_LOOP_for_for_for_asn_4996});
  assign buf_acc_data_4_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4986 , CONVOLUTION_LOOP_for_for_for_asn_4988
      , CONVOLUTION_LOOP_for_for_for_asn_4990});
  assign buf_acc_data_4_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4980 , CONVOLUTION_LOOP_for_for_for_asn_4982
      , CONVOLUTION_LOOP_for_for_for_asn_4984});
  assign buf_acc_data_4_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_4_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4974 , CONVOLUTION_LOOP_for_for_for_asn_4976
      , CONVOLUTION_LOOP_for_for_for_asn_4978});
  assign buf_acc_data_5_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4968 , CONVOLUTION_LOOP_for_for_for_asn_4970
      , CONVOLUTION_LOOP_for_for_for_asn_4972});
  assign buf_acc_data_5_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4962 , CONVOLUTION_LOOP_for_for_for_asn_4964
      , CONVOLUTION_LOOP_for_for_for_asn_4966});
  assign buf_acc_data_5_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4956 , CONVOLUTION_LOOP_for_for_for_asn_4958
      , CONVOLUTION_LOOP_for_for_for_asn_4960});
  assign buf_acc_data_5_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4950 , CONVOLUTION_LOOP_for_for_for_asn_4952
      , CONVOLUTION_LOOP_for_for_for_asn_4954});
  assign buf_acc_data_5_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4944 , CONVOLUTION_LOOP_for_for_for_asn_4946
      , CONVOLUTION_LOOP_for_for_for_asn_4948});
  assign buf_acc_data_5_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4938 , CONVOLUTION_LOOP_for_for_for_asn_4940
      , CONVOLUTION_LOOP_for_for_for_asn_4942});
  assign buf_acc_data_5_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4932 , CONVOLUTION_LOOP_for_for_for_asn_4934
      , CONVOLUTION_LOOP_for_for_for_asn_4936});
  assign buf_acc_data_5_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4926 , CONVOLUTION_LOOP_for_for_for_asn_4928
      , CONVOLUTION_LOOP_for_for_for_asn_4930});
  assign buf_acc_data_5_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4920 , CONVOLUTION_LOOP_for_for_for_asn_4922
      , CONVOLUTION_LOOP_for_for_for_asn_4924});
  assign buf_acc_data_5_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4914 , CONVOLUTION_LOOP_for_for_for_asn_4916
      , CONVOLUTION_LOOP_for_for_for_asn_4918});
  assign buf_acc_data_5_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4908 , CONVOLUTION_LOOP_for_for_for_asn_4910
      , CONVOLUTION_LOOP_for_for_for_asn_4912});
  assign buf_acc_data_5_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4902 , CONVOLUTION_LOOP_for_for_for_asn_4904
      , CONVOLUTION_LOOP_for_for_for_asn_4906});
  assign buf_acc_data_5_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4896 , CONVOLUTION_LOOP_for_for_for_asn_4898
      , CONVOLUTION_LOOP_for_for_for_asn_4900});
  assign buf_acc_data_5_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4890 , CONVOLUTION_LOOP_for_for_for_asn_4892
      , CONVOLUTION_LOOP_for_for_for_asn_4894});
  assign buf_acc_data_5_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4884 , CONVOLUTION_LOOP_for_for_for_asn_4886
      , CONVOLUTION_LOOP_for_for_for_asn_4888});
  assign buf_acc_data_5_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4878 , CONVOLUTION_LOOP_for_for_for_asn_4880
      , CONVOLUTION_LOOP_for_for_for_asn_4882});
  assign buf_acc_data_5_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4872 , CONVOLUTION_LOOP_for_for_for_asn_4874
      , CONVOLUTION_LOOP_for_for_for_asn_4876});
  assign buf_acc_data_5_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_5_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4866 , CONVOLUTION_LOOP_for_for_for_asn_4868
      , CONVOLUTION_LOOP_for_for_for_asn_4870});
  assign buf_acc_data_6_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4860 , CONVOLUTION_LOOP_for_for_for_asn_4862
      , CONVOLUTION_LOOP_for_for_for_asn_4864});
  assign buf_acc_data_6_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4854 , CONVOLUTION_LOOP_for_for_for_asn_4856
      , CONVOLUTION_LOOP_for_for_for_asn_4858});
  assign buf_acc_data_6_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4848 , CONVOLUTION_LOOP_for_for_for_asn_4850
      , CONVOLUTION_LOOP_for_for_for_asn_4852});
  assign buf_acc_data_6_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4842 , CONVOLUTION_LOOP_for_for_for_asn_4844
      , CONVOLUTION_LOOP_for_for_for_asn_4846});
  assign buf_acc_data_6_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4836 , CONVOLUTION_LOOP_for_for_for_asn_4838
      , CONVOLUTION_LOOP_for_for_for_asn_4840});
  assign buf_acc_data_6_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4830 , CONVOLUTION_LOOP_for_for_for_asn_4832
      , CONVOLUTION_LOOP_for_for_for_asn_4834});
  assign buf_acc_data_6_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4824 , CONVOLUTION_LOOP_for_for_for_asn_4826
      , CONVOLUTION_LOOP_for_for_for_asn_4828});
  assign buf_acc_data_6_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4818 , CONVOLUTION_LOOP_for_for_for_asn_4820
      , CONVOLUTION_LOOP_for_for_for_asn_4822});
  assign buf_acc_data_6_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4812 , CONVOLUTION_LOOP_for_for_for_asn_4814
      , CONVOLUTION_LOOP_for_for_for_asn_4816});
  assign buf_acc_data_6_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4806 , CONVOLUTION_LOOP_for_for_for_asn_4808
      , CONVOLUTION_LOOP_for_for_for_asn_4810});
  assign buf_acc_data_6_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4800 , CONVOLUTION_LOOP_for_for_for_asn_4802
      , CONVOLUTION_LOOP_for_for_for_asn_4804});
  assign buf_acc_data_6_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4794 , CONVOLUTION_LOOP_for_for_for_asn_4796
      , CONVOLUTION_LOOP_for_for_for_asn_4798});
  assign buf_acc_data_6_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4788 , CONVOLUTION_LOOP_for_for_for_asn_4790
      , CONVOLUTION_LOOP_for_for_for_asn_4792});
  assign buf_acc_data_6_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4782 , CONVOLUTION_LOOP_for_for_for_asn_4784
      , CONVOLUTION_LOOP_for_for_for_asn_4786});
  assign buf_acc_data_6_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4776 , CONVOLUTION_LOOP_for_for_for_asn_4778
      , CONVOLUTION_LOOP_for_for_for_asn_4780});
  assign buf_acc_data_6_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4770 , CONVOLUTION_LOOP_for_for_for_asn_4772
      , CONVOLUTION_LOOP_for_for_for_asn_4774});
  assign buf_acc_data_6_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4764 , CONVOLUTION_LOOP_for_for_for_asn_4766
      , CONVOLUTION_LOOP_for_for_for_asn_4768});
  assign buf_acc_data_6_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_6_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4758 , CONVOLUTION_LOOP_for_for_for_asn_4760
      , CONVOLUTION_LOOP_for_for_for_asn_4762});
  assign buf_acc_data_7_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4752 , CONVOLUTION_LOOP_for_for_for_asn_4754
      , CONVOLUTION_LOOP_for_for_for_asn_4756});
  assign buf_acc_data_7_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4746 , CONVOLUTION_LOOP_for_for_for_asn_4748
      , CONVOLUTION_LOOP_for_for_for_asn_4750});
  assign buf_acc_data_7_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4740 , CONVOLUTION_LOOP_for_for_for_asn_4742
      , CONVOLUTION_LOOP_for_for_for_asn_4744});
  assign buf_acc_data_7_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4734 , CONVOLUTION_LOOP_for_for_for_asn_4736
      , CONVOLUTION_LOOP_for_for_for_asn_4738});
  assign buf_acc_data_7_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4728 , CONVOLUTION_LOOP_for_for_for_asn_4730
      , CONVOLUTION_LOOP_for_for_for_asn_4732});
  assign buf_acc_data_7_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4722 , CONVOLUTION_LOOP_for_for_for_asn_4724
      , CONVOLUTION_LOOP_for_for_for_asn_4726});
  assign buf_acc_data_7_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4716 , CONVOLUTION_LOOP_for_for_for_asn_4718
      , CONVOLUTION_LOOP_for_for_for_asn_4720});
  assign buf_acc_data_7_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4710 , CONVOLUTION_LOOP_for_for_for_asn_4712
      , CONVOLUTION_LOOP_for_for_for_asn_4714});
  assign buf_acc_data_7_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4704 , CONVOLUTION_LOOP_for_for_for_asn_4706
      , CONVOLUTION_LOOP_for_for_for_asn_4708});
  assign buf_acc_data_7_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4698 , CONVOLUTION_LOOP_for_for_for_asn_4700
      , CONVOLUTION_LOOP_for_for_for_asn_4702});
  assign buf_acc_data_7_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4692 , CONVOLUTION_LOOP_for_for_for_asn_4694
      , CONVOLUTION_LOOP_for_for_for_asn_4696});
  assign buf_acc_data_7_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4686 , CONVOLUTION_LOOP_for_for_for_asn_4688
      , CONVOLUTION_LOOP_for_for_for_asn_4690});
  assign buf_acc_data_7_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4680 , CONVOLUTION_LOOP_for_for_for_asn_4682
      , CONVOLUTION_LOOP_for_for_for_asn_4684});
  assign buf_acc_data_7_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4674 , CONVOLUTION_LOOP_for_for_for_asn_4676
      , CONVOLUTION_LOOP_for_for_for_asn_4678});
  assign buf_acc_data_7_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4668 , CONVOLUTION_LOOP_for_for_for_asn_4670
      , CONVOLUTION_LOOP_for_for_for_asn_4672});
  assign buf_acc_data_7_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4662 , CONVOLUTION_LOOP_for_for_for_asn_4664
      , CONVOLUTION_LOOP_for_for_for_asn_4666});
  assign buf_acc_data_7_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4656 , CONVOLUTION_LOOP_for_for_for_asn_4658
      , CONVOLUTION_LOOP_for_for_for_asn_4660});
  assign buf_acc_data_7_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_7_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4650 , CONVOLUTION_LOOP_for_for_for_asn_4652
      , CONVOLUTION_LOOP_for_for_for_asn_4654});
  assign buf_acc_data_8_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4644 , CONVOLUTION_LOOP_for_for_for_asn_4646
      , CONVOLUTION_LOOP_for_for_for_asn_4648});
  assign buf_acc_data_8_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4638 , CONVOLUTION_LOOP_for_for_for_asn_4640
      , CONVOLUTION_LOOP_for_for_for_asn_4642});
  assign buf_acc_data_8_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4632 , CONVOLUTION_LOOP_for_for_for_asn_4634
      , CONVOLUTION_LOOP_for_for_for_asn_4636});
  assign buf_acc_data_8_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4626 , CONVOLUTION_LOOP_for_for_for_asn_4628
      , CONVOLUTION_LOOP_for_for_for_asn_4630});
  assign buf_acc_data_8_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4620 , CONVOLUTION_LOOP_for_for_for_asn_4622
      , CONVOLUTION_LOOP_for_for_for_asn_4624});
  assign buf_acc_data_8_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4614 , CONVOLUTION_LOOP_for_for_for_asn_4616
      , CONVOLUTION_LOOP_for_for_for_asn_4618});
  assign buf_acc_data_8_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4608 , CONVOLUTION_LOOP_for_for_for_asn_4610
      , CONVOLUTION_LOOP_for_for_for_asn_4612});
  assign buf_acc_data_8_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4602 , CONVOLUTION_LOOP_for_for_for_asn_4604
      , CONVOLUTION_LOOP_for_for_for_asn_4606});
  assign buf_acc_data_8_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4596 , CONVOLUTION_LOOP_for_for_for_asn_4598
      , CONVOLUTION_LOOP_for_for_for_asn_4600});
  assign buf_acc_data_8_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4590 , CONVOLUTION_LOOP_for_for_for_asn_4592
      , CONVOLUTION_LOOP_for_for_for_asn_4594});
  assign buf_acc_data_8_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4584 , CONVOLUTION_LOOP_for_for_for_asn_4586
      , CONVOLUTION_LOOP_for_for_for_asn_4588});
  assign buf_acc_data_8_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4578 , CONVOLUTION_LOOP_for_for_for_asn_4580
      , CONVOLUTION_LOOP_for_for_for_asn_4582});
  assign buf_acc_data_8_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4572 , CONVOLUTION_LOOP_for_for_for_asn_4574
      , CONVOLUTION_LOOP_for_for_for_asn_4576});
  assign buf_acc_data_8_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4566 , CONVOLUTION_LOOP_for_for_for_asn_4568
      , CONVOLUTION_LOOP_for_for_for_asn_4570});
  assign buf_acc_data_8_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4560 , CONVOLUTION_LOOP_for_for_for_asn_4562
      , CONVOLUTION_LOOP_for_for_for_asn_4564});
  assign buf_acc_data_8_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4554 , CONVOLUTION_LOOP_for_for_for_asn_4556
      , CONVOLUTION_LOOP_for_for_for_asn_4558});
  assign buf_acc_data_8_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4548 , CONVOLUTION_LOOP_for_for_for_asn_4550
      , CONVOLUTION_LOOP_for_for_for_asn_4552});
  assign buf_acc_data_8_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_8_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4542 , CONVOLUTION_LOOP_for_for_for_asn_4544
      , CONVOLUTION_LOOP_for_for_for_asn_4546});
  assign buf_acc_data_9_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4536 , CONVOLUTION_LOOP_for_for_for_asn_4538
      , CONVOLUTION_LOOP_for_for_for_asn_4540});
  assign buf_acc_data_9_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4530 , CONVOLUTION_LOOP_for_for_for_asn_4532
      , CONVOLUTION_LOOP_for_for_for_asn_4534});
  assign buf_acc_data_9_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4524 , CONVOLUTION_LOOP_for_for_for_asn_4526
      , CONVOLUTION_LOOP_for_for_for_asn_4528});
  assign buf_acc_data_9_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4518 , CONVOLUTION_LOOP_for_for_for_asn_4520
      , CONVOLUTION_LOOP_for_for_for_asn_4522});
  assign buf_acc_data_9_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4512 , CONVOLUTION_LOOP_for_for_for_asn_4514
      , CONVOLUTION_LOOP_for_for_for_asn_4516});
  assign buf_acc_data_9_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4506 , CONVOLUTION_LOOP_for_for_for_asn_4508
      , CONVOLUTION_LOOP_for_for_for_asn_4510});
  assign buf_acc_data_9_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4500 , CONVOLUTION_LOOP_for_for_for_asn_4502
      , CONVOLUTION_LOOP_for_for_for_asn_4504});
  assign buf_acc_data_9_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4494 , CONVOLUTION_LOOP_for_for_for_asn_4496
      , CONVOLUTION_LOOP_for_for_for_asn_4498});
  assign buf_acc_data_9_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4488 , CONVOLUTION_LOOP_for_for_for_asn_4490
      , CONVOLUTION_LOOP_for_for_for_asn_4492});
  assign buf_acc_data_9_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4482 , CONVOLUTION_LOOP_for_for_for_asn_4484
      , CONVOLUTION_LOOP_for_for_for_asn_4486});
  assign buf_acc_data_9_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4476 , CONVOLUTION_LOOP_for_for_for_asn_4478
      , CONVOLUTION_LOOP_for_for_for_asn_4480});
  assign buf_acc_data_9_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4470 , CONVOLUTION_LOOP_for_for_for_asn_4472
      , CONVOLUTION_LOOP_for_for_for_asn_4474});
  assign buf_acc_data_9_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4464 , CONVOLUTION_LOOP_for_for_for_asn_4466
      , CONVOLUTION_LOOP_for_for_for_asn_4468});
  assign buf_acc_data_9_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4458 , CONVOLUTION_LOOP_for_for_for_asn_4460
      , CONVOLUTION_LOOP_for_for_for_asn_4462});
  assign buf_acc_data_9_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4452 , CONVOLUTION_LOOP_for_for_for_asn_4454
      , CONVOLUTION_LOOP_for_for_for_asn_4456});
  assign buf_acc_data_9_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4446 , CONVOLUTION_LOOP_for_for_for_asn_4448
      , CONVOLUTION_LOOP_for_for_for_asn_4450});
  assign buf_acc_data_9_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4440 , CONVOLUTION_LOOP_for_for_for_asn_4442
      , CONVOLUTION_LOOP_for_for_for_asn_4444});
  assign buf_acc_data_9_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_9_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4434 , CONVOLUTION_LOOP_for_for_for_asn_4436
      , CONVOLUTION_LOOP_for_for_for_asn_4438});
  assign buf_acc_data_10_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4428 , CONVOLUTION_LOOP_for_for_for_asn_4430
      , CONVOLUTION_LOOP_for_for_for_asn_4432});
  assign buf_acc_data_10_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4422 , CONVOLUTION_LOOP_for_for_for_asn_4424
      , CONVOLUTION_LOOP_for_for_for_asn_4426});
  assign buf_acc_data_10_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4416 , CONVOLUTION_LOOP_for_for_for_asn_4418
      , CONVOLUTION_LOOP_for_for_for_asn_4420});
  assign buf_acc_data_10_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4410 , CONVOLUTION_LOOP_for_for_for_asn_4412
      , CONVOLUTION_LOOP_for_for_for_asn_4414});
  assign buf_acc_data_10_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4404 , CONVOLUTION_LOOP_for_for_for_asn_4406
      , CONVOLUTION_LOOP_for_for_for_asn_4408});
  assign buf_acc_data_10_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4398 , CONVOLUTION_LOOP_for_for_for_asn_4400
      , CONVOLUTION_LOOP_for_for_for_asn_4402});
  assign buf_acc_data_10_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4392 , CONVOLUTION_LOOP_for_for_for_asn_4394
      , CONVOLUTION_LOOP_for_for_for_asn_4396});
  assign buf_acc_data_10_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4386 , CONVOLUTION_LOOP_for_for_for_asn_4388
      , CONVOLUTION_LOOP_for_for_for_asn_4390});
  assign buf_acc_data_10_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4380 , CONVOLUTION_LOOP_for_for_for_asn_4382
      , CONVOLUTION_LOOP_for_for_for_asn_4384});
  assign buf_acc_data_10_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4374 , CONVOLUTION_LOOP_for_for_for_asn_4376
      , CONVOLUTION_LOOP_for_for_for_asn_4378});
  assign buf_acc_data_10_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4368 , CONVOLUTION_LOOP_for_for_for_asn_4370
      , CONVOLUTION_LOOP_for_for_for_asn_4372});
  assign buf_acc_data_10_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4362 , CONVOLUTION_LOOP_for_for_for_asn_4364
      , CONVOLUTION_LOOP_for_for_for_asn_4366});
  assign buf_acc_data_10_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4356 , CONVOLUTION_LOOP_for_for_for_asn_4358
      , CONVOLUTION_LOOP_for_for_for_asn_4360});
  assign buf_acc_data_10_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4350 , CONVOLUTION_LOOP_for_for_for_asn_4352
      , CONVOLUTION_LOOP_for_for_for_asn_4354});
  assign buf_acc_data_10_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4344 , CONVOLUTION_LOOP_for_for_for_asn_4346
      , CONVOLUTION_LOOP_for_for_for_asn_4348});
  assign buf_acc_data_10_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4338 , CONVOLUTION_LOOP_for_for_for_asn_4340
      , CONVOLUTION_LOOP_for_for_for_asn_4342});
  assign buf_acc_data_10_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4332 , CONVOLUTION_LOOP_for_for_for_asn_4334
      , CONVOLUTION_LOOP_for_for_for_asn_4336});
  assign buf_acc_data_10_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_10_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4326 , CONVOLUTION_LOOP_for_for_for_asn_4328
      , CONVOLUTION_LOOP_for_for_for_asn_4330});
  assign buf_acc_data_11_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4320 , CONVOLUTION_LOOP_for_for_for_asn_4322
      , CONVOLUTION_LOOP_for_for_for_asn_4324});
  assign buf_acc_data_11_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4314 , CONVOLUTION_LOOP_for_for_for_asn_4316
      , CONVOLUTION_LOOP_for_for_for_asn_4318});
  assign buf_acc_data_11_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4308 , CONVOLUTION_LOOP_for_for_for_asn_4310
      , CONVOLUTION_LOOP_for_for_for_asn_4312});
  assign buf_acc_data_11_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4302 , CONVOLUTION_LOOP_for_for_for_asn_4304
      , CONVOLUTION_LOOP_for_for_for_asn_4306});
  assign buf_acc_data_11_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4296 , CONVOLUTION_LOOP_for_for_for_asn_4298
      , CONVOLUTION_LOOP_for_for_for_asn_4300});
  assign buf_acc_data_11_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4290 , CONVOLUTION_LOOP_for_for_for_asn_4292
      , CONVOLUTION_LOOP_for_for_for_asn_4294});
  assign buf_acc_data_11_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4284 , CONVOLUTION_LOOP_for_for_for_asn_4286
      , CONVOLUTION_LOOP_for_for_for_asn_4288});
  assign buf_acc_data_11_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4278 , CONVOLUTION_LOOP_for_for_for_asn_4280
      , CONVOLUTION_LOOP_for_for_for_asn_4282});
  assign buf_acc_data_11_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4272 , CONVOLUTION_LOOP_for_for_for_asn_4274
      , CONVOLUTION_LOOP_for_for_for_asn_4276});
  assign buf_acc_data_11_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4266 , CONVOLUTION_LOOP_for_for_for_asn_4268
      , CONVOLUTION_LOOP_for_for_for_asn_4270});
  assign buf_acc_data_11_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4260 , CONVOLUTION_LOOP_for_for_for_asn_4262
      , CONVOLUTION_LOOP_for_for_for_asn_4264});
  assign buf_acc_data_11_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4254 , CONVOLUTION_LOOP_for_for_for_asn_4256
      , CONVOLUTION_LOOP_for_for_for_asn_4258});
  assign buf_acc_data_11_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4248 , CONVOLUTION_LOOP_for_for_for_asn_4250
      , CONVOLUTION_LOOP_for_for_for_asn_4252});
  assign buf_acc_data_11_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4242 , CONVOLUTION_LOOP_for_for_for_asn_4244
      , CONVOLUTION_LOOP_for_for_for_asn_4246});
  assign buf_acc_data_11_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4236 , CONVOLUTION_LOOP_for_for_for_asn_4238
      , CONVOLUTION_LOOP_for_for_for_asn_4240});
  assign buf_acc_data_11_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4230 , CONVOLUTION_LOOP_for_for_for_asn_4232
      , CONVOLUTION_LOOP_for_for_for_asn_4234});
  assign buf_acc_data_11_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4224 , CONVOLUTION_LOOP_for_for_for_asn_4226
      , CONVOLUTION_LOOP_for_for_for_asn_4228});
  assign buf_acc_data_11_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_11_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4218 , CONVOLUTION_LOOP_for_for_for_asn_4220
      , CONVOLUTION_LOOP_for_for_for_asn_4222});
  assign buf_acc_data_12_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4212 , CONVOLUTION_LOOP_for_for_for_asn_4214
      , CONVOLUTION_LOOP_for_for_for_asn_4216});
  assign buf_acc_data_12_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4206 , CONVOLUTION_LOOP_for_for_for_asn_4208
      , CONVOLUTION_LOOP_for_for_for_asn_4210});
  assign buf_acc_data_12_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4200 , CONVOLUTION_LOOP_for_for_for_asn_4202
      , CONVOLUTION_LOOP_for_for_for_asn_4204});
  assign buf_acc_data_12_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4194 , CONVOLUTION_LOOP_for_for_for_asn_4196
      , CONVOLUTION_LOOP_for_for_for_asn_4198});
  assign buf_acc_data_12_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4188 , CONVOLUTION_LOOP_for_for_for_asn_4190
      , CONVOLUTION_LOOP_for_for_for_asn_4192});
  assign buf_acc_data_12_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4182 , CONVOLUTION_LOOP_for_for_for_asn_4184
      , CONVOLUTION_LOOP_for_for_for_asn_4186});
  assign buf_acc_data_12_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4176 , CONVOLUTION_LOOP_for_for_for_asn_4178
      , CONVOLUTION_LOOP_for_for_for_asn_4180});
  assign buf_acc_data_12_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4170 , CONVOLUTION_LOOP_for_for_for_asn_4172
      , CONVOLUTION_LOOP_for_for_for_asn_4174});
  assign buf_acc_data_12_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4164 , CONVOLUTION_LOOP_for_for_for_asn_4166
      , CONVOLUTION_LOOP_for_for_for_asn_4168});
  assign buf_acc_data_12_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4158 , CONVOLUTION_LOOP_for_for_for_asn_4160
      , CONVOLUTION_LOOP_for_for_for_asn_4162});
  assign buf_acc_data_12_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4152 , CONVOLUTION_LOOP_for_for_for_asn_4154
      , CONVOLUTION_LOOP_for_for_for_asn_4156});
  assign buf_acc_data_12_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4146 , CONVOLUTION_LOOP_for_for_for_asn_4148
      , CONVOLUTION_LOOP_for_for_for_asn_4150});
  assign buf_acc_data_12_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4140 , CONVOLUTION_LOOP_for_for_for_asn_4142
      , CONVOLUTION_LOOP_for_for_for_asn_4144});
  assign buf_acc_data_12_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4134 , CONVOLUTION_LOOP_for_for_for_asn_4136
      , CONVOLUTION_LOOP_for_for_for_asn_4138});
  assign buf_acc_data_12_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4128 , CONVOLUTION_LOOP_for_for_for_asn_4130
      , CONVOLUTION_LOOP_for_for_for_asn_4132});
  assign buf_acc_data_12_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4122 , CONVOLUTION_LOOP_for_for_for_asn_4124
      , CONVOLUTION_LOOP_for_for_for_asn_4126});
  assign buf_acc_data_12_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4116 , CONVOLUTION_LOOP_for_for_for_asn_4118
      , CONVOLUTION_LOOP_for_for_for_asn_4120});
  assign buf_acc_data_12_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_12_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4110 , CONVOLUTION_LOOP_for_for_for_asn_4112
      , CONVOLUTION_LOOP_for_for_for_asn_4114});
  assign buf_acc_data_13_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4104 , CONVOLUTION_LOOP_for_for_for_asn_4106
      , CONVOLUTION_LOOP_for_for_for_asn_4108});
  assign buf_acc_data_13_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4098 , CONVOLUTION_LOOP_for_for_for_asn_4100
      , CONVOLUTION_LOOP_for_for_for_asn_4102});
  assign buf_acc_data_13_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4092 , CONVOLUTION_LOOP_for_for_for_asn_4094
      , CONVOLUTION_LOOP_for_for_for_asn_4096});
  assign buf_acc_data_13_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4086 , CONVOLUTION_LOOP_for_for_for_asn_4088
      , CONVOLUTION_LOOP_for_for_for_asn_4090});
  assign buf_acc_data_13_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4080 , CONVOLUTION_LOOP_for_for_for_asn_4082
      , CONVOLUTION_LOOP_for_for_for_asn_4084});
  assign buf_acc_data_13_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4074 , CONVOLUTION_LOOP_for_for_for_asn_4076
      , CONVOLUTION_LOOP_for_for_for_asn_4078});
  assign buf_acc_data_13_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4068 , CONVOLUTION_LOOP_for_for_for_asn_4070
      , CONVOLUTION_LOOP_for_for_for_asn_4072});
  assign buf_acc_data_13_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4062 , CONVOLUTION_LOOP_for_for_for_asn_4064
      , CONVOLUTION_LOOP_for_for_for_asn_4066});
  assign buf_acc_data_13_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4056 , CONVOLUTION_LOOP_for_for_for_asn_4058
      , CONVOLUTION_LOOP_for_for_for_asn_4060});
  assign buf_acc_data_13_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4050 , CONVOLUTION_LOOP_for_for_for_asn_4052
      , CONVOLUTION_LOOP_for_for_for_asn_4054});
  assign buf_acc_data_13_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4044 , CONVOLUTION_LOOP_for_for_for_asn_4046
      , CONVOLUTION_LOOP_for_for_for_asn_4048});
  assign buf_acc_data_13_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4038 , CONVOLUTION_LOOP_for_for_for_asn_4040
      , CONVOLUTION_LOOP_for_for_for_asn_4042});
  assign buf_acc_data_13_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4032 , CONVOLUTION_LOOP_for_for_for_asn_4034
      , CONVOLUTION_LOOP_for_for_for_asn_4036});
  assign buf_acc_data_13_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4026 , CONVOLUTION_LOOP_for_for_for_asn_4028
      , CONVOLUTION_LOOP_for_for_for_asn_4030});
  assign buf_acc_data_13_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4020 , CONVOLUTION_LOOP_for_for_for_asn_4022
      , CONVOLUTION_LOOP_for_for_for_asn_4024});
  assign buf_acc_data_13_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4014 , CONVOLUTION_LOOP_for_for_for_asn_4016
      , CONVOLUTION_LOOP_for_for_for_asn_4018});
  assign buf_acc_data_13_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4008 , CONVOLUTION_LOOP_for_for_for_asn_4010
      , CONVOLUTION_LOOP_for_for_for_asn_4012});
  assign buf_acc_data_13_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_13_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4002 , CONVOLUTION_LOOP_for_for_for_asn_4004
      , CONVOLUTION_LOOP_for_for_for_asn_4006});
  assign buf_acc_data_14_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3996 , CONVOLUTION_LOOP_for_for_for_asn_3998
      , CONVOLUTION_LOOP_for_for_for_asn_4000});
  assign buf_acc_data_14_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3990 , CONVOLUTION_LOOP_for_for_for_asn_3992
      , CONVOLUTION_LOOP_for_for_for_asn_3994});
  assign buf_acc_data_14_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3984 , CONVOLUTION_LOOP_for_for_for_asn_3986
      , CONVOLUTION_LOOP_for_for_for_asn_3988});
  assign buf_acc_data_14_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3978 , CONVOLUTION_LOOP_for_for_for_asn_3980
      , CONVOLUTION_LOOP_for_for_for_asn_3982});
  assign buf_acc_data_14_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3972 , CONVOLUTION_LOOP_for_for_for_asn_3974
      , CONVOLUTION_LOOP_for_for_for_asn_3976});
  assign buf_acc_data_14_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3966 , CONVOLUTION_LOOP_for_for_for_asn_3968
      , CONVOLUTION_LOOP_for_for_for_asn_3970});
  assign buf_acc_data_14_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3960 , CONVOLUTION_LOOP_for_for_for_asn_3962
      , CONVOLUTION_LOOP_for_for_for_asn_3964});
  assign buf_acc_data_14_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3954 , CONVOLUTION_LOOP_for_for_for_asn_3956
      , CONVOLUTION_LOOP_for_for_for_asn_3958});
  assign buf_acc_data_14_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3948 , CONVOLUTION_LOOP_for_for_for_asn_3950
      , CONVOLUTION_LOOP_for_for_for_asn_3952});
  assign buf_acc_data_14_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3942 , CONVOLUTION_LOOP_for_for_for_asn_3944
      , CONVOLUTION_LOOP_for_for_for_asn_3946});
  assign buf_acc_data_14_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3936 , CONVOLUTION_LOOP_for_for_for_asn_3938
      , CONVOLUTION_LOOP_for_for_for_asn_3940});
  assign buf_acc_data_14_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3930 , CONVOLUTION_LOOP_for_for_for_asn_3932
      , CONVOLUTION_LOOP_for_for_for_asn_3934});
  assign buf_acc_data_14_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3924 , CONVOLUTION_LOOP_for_for_for_asn_3926
      , CONVOLUTION_LOOP_for_for_for_asn_3928});
  assign buf_acc_data_14_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3918 , CONVOLUTION_LOOP_for_for_for_asn_3920
      , CONVOLUTION_LOOP_for_for_for_asn_3922});
  assign buf_acc_data_14_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3912 , CONVOLUTION_LOOP_for_for_for_asn_3914
      , CONVOLUTION_LOOP_for_for_for_asn_3916});
  assign buf_acc_data_14_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3906 , CONVOLUTION_LOOP_for_for_for_asn_3908
      , CONVOLUTION_LOOP_for_for_for_asn_3910});
  assign buf_acc_data_14_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3900 , CONVOLUTION_LOOP_for_for_for_asn_3902
      , CONVOLUTION_LOOP_for_for_for_asn_3904});
  assign buf_acc_data_14_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_14_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3894 , CONVOLUTION_LOOP_for_for_for_asn_3896
      , CONVOLUTION_LOOP_for_for_for_asn_3898});
  assign buf_acc_data_15_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3888 , CONVOLUTION_LOOP_for_for_for_asn_3890
      , CONVOLUTION_LOOP_for_for_for_asn_3892});
  assign buf_acc_data_15_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3882 , CONVOLUTION_LOOP_for_for_for_asn_3884
      , CONVOLUTION_LOOP_for_for_for_asn_3886});
  assign buf_acc_data_15_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3876 , CONVOLUTION_LOOP_for_for_for_asn_3878
      , CONVOLUTION_LOOP_for_for_for_asn_3880});
  assign buf_acc_data_15_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3870 , CONVOLUTION_LOOP_for_for_for_asn_3872
      , CONVOLUTION_LOOP_for_for_for_asn_3874});
  assign buf_acc_data_15_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3864 , CONVOLUTION_LOOP_for_for_for_asn_3866
      , CONVOLUTION_LOOP_for_for_for_asn_3868});
  assign buf_acc_data_15_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3858 , CONVOLUTION_LOOP_for_for_for_asn_3860
      , CONVOLUTION_LOOP_for_for_for_asn_3862});
  assign buf_acc_data_15_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3852 , CONVOLUTION_LOOP_for_for_for_asn_3854
      , CONVOLUTION_LOOP_for_for_for_asn_3856});
  assign buf_acc_data_15_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3846 , CONVOLUTION_LOOP_for_for_for_asn_3848
      , CONVOLUTION_LOOP_for_for_for_asn_3850});
  assign buf_acc_data_15_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3840 , CONVOLUTION_LOOP_for_for_for_asn_3842
      , CONVOLUTION_LOOP_for_for_for_asn_3844});
  assign buf_acc_data_15_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3834 , CONVOLUTION_LOOP_for_for_for_asn_3836
      , CONVOLUTION_LOOP_for_for_for_asn_3838});
  assign buf_acc_data_15_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3828 , CONVOLUTION_LOOP_for_for_for_asn_3830
      , CONVOLUTION_LOOP_for_for_for_asn_3832});
  assign buf_acc_data_15_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3822 , CONVOLUTION_LOOP_for_for_for_asn_3824
      , CONVOLUTION_LOOP_for_for_for_asn_3826});
  assign buf_acc_data_15_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3816 , CONVOLUTION_LOOP_for_for_for_asn_3818
      , CONVOLUTION_LOOP_for_for_for_asn_3820});
  assign buf_acc_data_15_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3810 , CONVOLUTION_LOOP_for_for_for_asn_3812
      , CONVOLUTION_LOOP_for_for_for_asn_3814});
  assign buf_acc_data_15_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3804 , CONVOLUTION_LOOP_for_for_for_asn_3806
      , CONVOLUTION_LOOP_for_for_for_asn_3808});
  assign buf_acc_data_15_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3798 , CONVOLUTION_LOOP_for_for_for_asn_3800
      , CONVOLUTION_LOOP_for_for_for_asn_3802});
  assign buf_acc_data_15_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3792 , CONVOLUTION_LOOP_for_for_for_asn_3794
      , CONVOLUTION_LOOP_for_for_for_asn_3796});
  assign buf_acc_data_15_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_15_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3786 , CONVOLUTION_LOOP_for_for_for_asn_3788
      , CONVOLUTION_LOOP_for_for_for_asn_3790});
  assign buf_acc_data_16_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3780 , CONVOLUTION_LOOP_for_for_for_asn_3782
      , CONVOLUTION_LOOP_for_for_for_asn_3784});
  assign buf_acc_data_16_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3774 , CONVOLUTION_LOOP_for_for_for_asn_3776
      , CONVOLUTION_LOOP_for_for_for_asn_3778});
  assign buf_acc_data_16_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3768 , CONVOLUTION_LOOP_for_for_for_asn_3770
      , CONVOLUTION_LOOP_for_for_for_asn_3772});
  assign buf_acc_data_16_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3762 , CONVOLUTION_LOOP_for_for_for_asn_3764
      , CONVOLUTION_LOOP_for_for_for_asn_3766});
  assign buf_acc_data_16_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3756 , CONVOLUTION_LOOP_for_for_for_asn_3758
      , CONVOLUTION_LOOP_for_for_for_asn_3760});
  assign buf_acc_data_16_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3750 , CONVOLUTION_LOOP_for_for_for_asn_3752
      , CONVOLUTION_LOOP_for_for_for_asn_3754});
  assign buf_acc_data_16_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3744 , CONVOLUTION_LOOP_for_for_for_asn_3746
      , CONVOLUTION_LOOP_for_for_for_asn_3748});
  assign buf_acc_data_16_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3738 , CONVOLUTION_LOOP_for_for_for_asn_3740
      , CONVOLUTION_LOOP_for_for_for_asn_3742});
  assign buf_acc_data_16_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3732 , CONVOLUTION_LOOP_for_for_for_asn_3734
      , CONVOLUTION_LOOP_for_for_for_asn_3736});
  assign buf_acc_data_16_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3726 , CONVOLUTION_LOOP_for_for_for_asn_3728
      , CONVOLUTION_LOOP_for_for_for_asn_3730});
  assign buf_acc_data_16_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3720 , CONVOLUTION_LOOP_for_for_for_asn_3722
      , CONVOLUTION_LOOP_for_for_for_asn_3724});
  assign buf_acc_data_16_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3714 , CONVOLUTION_LOOP_for_for_for_asn_3716
      , CONVOLUTION_LOOP_for_for_for_asn_3718});
  assign buf_acc_data_16_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3708 , CONVOLUTION_LOOP_for_for_for_asn_3710
      , CONVOLUTION_LOOP_for_for_for_asn_3712});
  assign buf_acc_data_16_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3702 , CONVOLUTION_LOOP_for_for_for_asn_3704
      , CONVOLUTION_LOOP_for_for_for_asn_3706});
  assign buf_acc_data_16_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3696 , CONVOLUTION_LOOP_for_for_for_asn_3698
      , CONVOLUTION_LOOP_for_for_for_asn_3700});
  assign buf_acc_data_16_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3690 , CONVOLUTION_LOOP_for_for_for_asn_3692
      , CONVOLUTION_LOOP_for_for_for_asn_3694});
  assign buf_acc_data_16_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3684 , CONVOLUTION_LOOP_for_for_for_asn_3686
      , CONVOLUTION_LOOP_for_for_for_asn_3688});
  assign buf_acc_data_16_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_16_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3678 , CONVOLUTION_LOOP_for_for_for_asn_3680
      , CONVOLUTION_LOOP_for_for_for_asn_3682});
  assign buf_acc_data_17_0_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_0_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3672 , CONVOLUTION_LOOP_for_for_for_asn_3674
      , CONVOLUTION_LOOP_for_for_for_asn_3676});
  assign buf_acc_data_17_1_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_1_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3666 , CONVOLUTION_LOOP_for_for_for_asn_3668
      , CONVOLUTION_LOOP_for_for_for_asn_3670});
  assign buf_acc_data_17_2_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_2_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3660 , CONVOLUTION_LOOP_for_for_for_asn_3662
      , CONVOLUTION_LOOP_for_for_for_asn_3664});
  assign buf_acc_data_17_3_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_3_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3654 , CONVOLUTION_LOOP_for_for_for_asn_3656
      , CONVOLUTION_LOOP_for_for_for_asn_3658});
  assign buf_acc_data_17_4_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_4_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3648 , CONVOLUTION_LOOP_for_for_for_asn_3650
      , CONVOLUTION_LOOP_for_for_for_asn_3652});
  assign buf_acc_data_17_5_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_5_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3642 , CONVOLUTION_LOOP_for_for_for_asn_3644
      , CONVOLUTION_LOOP_for_for_for_asn_3646});
  assign buf_acc_data_17_6_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_6_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3636 , CONVOLUTION_LOOP_for_for_for_asn_3638
      , CONVOLUTION_LOOP_for_for_for_asn_3640});
  assign buf_acc_data_17_7_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_7_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3630 , CONVOLUTION_LOOP_for_for_for_asn_3632
      , CONVOLUTION_LOOP_for_for_for_asn_3634});
  assign buf_acc_data_17_8_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_8_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3624 , CONVOLUTION_LOOP_for_for_for_asn_3626
      , CONVOLUTION_LOOP_for_for_for_asn_3628});
  assign buf_acc_data_17_9_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_9_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3618 , CONVOLUTION_LOOP_for_for_for_asn_3620
      , CONVOLUTION_LOOP_for_for_for_asn_3622});
  assign buf_acc_data_17_10_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_10_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3612 , CONVOLUTION_LOOP_for_for_for_asn_3614
      , CONVOLUTION_LOOP_for_for_for_asn_3616});
  assign buf_acc_data_17_11_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_11_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3606 , CONVOLUTION_LOOP_for_for_for_asn_3608
      , CONVOLUTION_LOOP_for_for_for_asn_3610});
  assign buf_acc_data_17_12_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_12_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3600 , CONVOLUTION_LOOP_for_for_for_asn_3602
      , CONVOLUTION_LOOP_for_for_for_asn_3604});
  assign buf_acc_data_17_13_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_13_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3594 , CONVOLUTION_LOOP_for_for_for_asn_3596
      , CONVOLUTION_LOOP_for_for_for_asn_3598});
  assign buf_acc_data_17_14_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_14_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3588 , CONVOLUTION_LOOP_for_for_for_asn_3590
      , CONVOLUTION_LOOP_for_for_for_asn_3592});
  assign buf_acc_data_17_15_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_15_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3582 , CONVOLUTION_LOOP_for_for_for_asn_3584
      , CONVOLUTION_LOOP_for_for_for_asn_3586});
  assign buf_acc_data_17_16_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_16_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3576 , CONVOLUTION_LOOP_for_for_for_asn_3578
      , CONVOLUTION_LOOP_for_for_for_asn_3580});
  assign buf_acc_data_17_17_45_1_sva_dfm_1 = MUX1HOT_v_45_3_2(buf_acc_data_17_17_45_1_sva,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3570 , CONVOLUTION_LOOP_for_for_for_asn_3572
      , CONVOLUTION_LOOP_for_for_for_asn_3574});
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_nl = (z_out_7[15]) & ((z_out_7[14:0]!=15'b000000000000000)
      | (CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1[0]));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1 = CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1
      + conv_u2s_1_49(CONVOLUTION_LOOP_for_for_for_for_for_and_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[48:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[48])
      & (~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[47:46]==2'b11)));
  assign CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[48])
      | (~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[47:46]!=2'b00))));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1 = conv_s2u_47_49({CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
      , CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
      , CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1})
      + conv_s2u_48_49(z_out_7[63:16]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1[48:0];
  assign LOAD_LOOP_LOAD_LOOP_if_and_tmp = (LOAD_LOOP_i_lpi_2_mx1 == (operator_32_false_acc_psp_sva_1[15:0]))
      & (operator_32_false_acc_psp_sva_1[32:16]==17'b00000000000000000);
  assign nl_operator_32_false_acc_psp_sva_1 = conv_u2s_32_33(z_out_10) + 33'b111111111111111111111111111111111;
  assign operator_32_false_acc_psp_sva_1 = nl_operator_32_false_acc_psp_sva_1[32:0];
  assign nl_PADDING_LOOP_for_for_aelse_1_acc_1_nl = conv_u2u_8_9({(~ n_h_in_acc_psp_sva)
      , (~ (conf_info_crt_sva_231_0[160]))}) + conv_u2u_8_9(pad_sva) + 9'b000000001;
  assign PADDING_LOOP_for_for_aelse_1_acc_1_nl = nl_PADDING_LOOP_for_for_aelse_1_acc_1_nl[8:0];
  assign nl_PADDING_LOOP_for_for_aelse_1_acc_nl = conv_u2u_9_10(PADDING_LOOP_for_for_aelse_1_acc_1_nl)
      + conv_s2u_9_10({4'b1000 , PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5});
  assign PADDING_LOOP_for_for_aelse_1_acc_nl = nl_PADDING_LOOP_for_for_aelse_1_acc_nl[9:0];
  assign PADDING_LOOP_for_for_aelse_1_acc_itm_9_1 = readslicef_10_1_9(PADDING_LOOP_for_for_aelse_1_acc_nl);
  assign PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5 = MUX_v_5_2_2(5'b00000, PADDING_LOOP_for_for_col_4_0_lpi_2,
      lfst_exit_PADDING_LOOP_for_lpi_2);
  assign exit_PADDING_LOOP_sva_2 = ~((~((PADDING_LOOP_chan_5_0_lpi_2_4_0 == (z_out_4[4:0]))
      & CONVOLUTION_LOOP_for_if_nor_cse)) | (z_out_4[8]));
  assign nl_operator_8_false_2_acc_nl = conv_u2s_4_5(PADDING_LOOP_for_row_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_2_acc_nl = nl_operator_8_false_2_acc_nl[4:0];
  assign operator_8_false_2_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_2_acc_nl);
  assign nl_PADDING_LOOP_for_row_4_0_sva_2 = PADDING_LOOP_for_row_4_0_lpi_2 + 5'b00001;
  assign PADDING_LOOP_for_row_4_0_sva_2 = nl_PADDING_LOOP_for_row_4_0_sva_2[4:0];
  assign PADDING_LOOP_for_if_equal_tmp = PADDING_LOOP_for_row_4_0_lpi_2 == (operator_8_false_2_acc_tmp[4:0]);
  assign exit_PADDING_LOOP_for_sva_5 = ~((~(PADDING_LOOP_for_if_equal_tmp & (operator_8_false_2_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_2_acc_tmp[8]));
  assign nl_operator_8_false_2_acc_tmp = conv_u2s_8_9({n_w_in_acc_psp_sva , (conf_info_crt_sva_231_0[192])})
      + 9'b111111111;
  assign operator_8_false_2_acc_tmp = nl_operator_8_false_2_acc_tmp[8:0];
  assign nl_operator_8_false_3_acc_nl = conv_u2s_4_5(PADDING_LOOP_for_for_col_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_3_acc_nl = nl_operator_8_false_3_acc_nl[4:0];
  assign operator_8_false_3_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_3_acc_nl);
  assign nl_PADDING_LOOP_for_for_col_4_0_sva_2 = PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5
      + 5'b00001;
  assign PADDING_LOOP_for_for_col_4_0_sva_2 = nl_PADDING_LOOP_for_for_col_4_0_sva_2[4:0];
  assign PADDING_LOOP_for_mux_1_nl = MUX_s_1_2_2(exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0,
      exit_PADDING_LOOP_for_lpi_2_dfm_1, and_dcpl_79);
  assign exit_PADDING_LOOP_for_lpi_2_dfm_4 = PADDING_LOOP_for_mux_1_nl & exit_PADDING_LOOP_for_for_lpi_2_dfm_1;
  assign exit_PADDING_LOOP_for_for_lpi_2_dfm_1 = ~(operator_8_false_3_acc_itm_4_1
      & ((~(PADDING_LOOP_for_for_if_1_equal_tmp & (operator_8_false_1_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_1_acc_tmp[8])));
  assign PADDING_LOOP_for_for_if_1_equal_tmp = PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5
      == (operator_8_false_1_acc_tmp[4:0]);
  assign nl_operator_8_false_1_acc_tmp = conv_u2s_8_9({n_h_in_acc_psp_sva , (conf_info_crt_sva_231_0[160])})
      + 9'b111111111;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[8:0];
  assign nl_CONVOLUTION_LOOP_acc_tmp = conv_u2u_5_6(CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0)
      + 6'b000001;
  assign CONVOLUTION_LOOP_acc_tmp = nl_CONVOLUTION_LOOP_acc_tmp[5:0];
  assign CONVOLUTION_LOOP_if_equal_tmp = CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0 == (operator_8_false_10_acc_tmp[4:0]);
  assign exit_CONVOLUTION_LOOP_sva_2 = ~((~(CONVOLUTION_LOOP_if_equal_tmp & (operator_8_false_10_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_10_acc_tmp[8]));
  assign nl_operator_8_false_10_acc_tmp = conv_u2s_8_9(conf_info_crt_sva_231_0[71:64])
      + 9'b111111111;
  assign operator_8_false_10_acc_tmp = nl_operator_8_false_10_acc_tmp[8:0];
  assign nl_CONVOLUTION_LOOP_for_acc_tmp = conv_u2u_5_6(CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1)
      + 6'b000001;
  assign CONVOLUTION_LOOP_for_acc_tmp = nl_CONVOLUTION_LOOP_for_acc_tmp[5:0];
  assign CONVOLUTION_LOOP_for_if_nor_cse = ~((z_out_4[7:5]!=3'b000));
  assign nl_operator_8_false_6_acc_nl = conv_u2s_4_5(CONVOLUTION_LOOP_for_for_i_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_6_acc_nl = nl_operator_8_false_6_acc_nl[4:0];
  assign operator_8_false_6_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_6_acc_nl);
  assign nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2 = CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6
      + 5'b00001;
  assign CONVOLUTION_LOOP_for_for_i_4_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2[4:0];
  assign CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6 = MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_for_i_4_0_lpi_2,
      lfst_exit_CONVOLUTION_LOOP_for_lpi_2);
  assign CONVOLUTION_LOOP_for_for_if_equal_tmp = CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6
      == (operator_8_false_8_acc_tmp[4:0]);
  assign nl_operator_8_false_8_acc_tmp = conv_u2s_8_9(n_w_out_lpi_1_dfm) + 9'b111111111;
  assign operator_8_false_8_acc_tmp = nl_operator_8_false_8_acc_tmp[8:0];
  assign nl_operator_8_false_7_acc_nl = conv_u2s_4_5(CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_7_acc_nl = nl_operator_8_false_7_acc_nl[4:0];
  assign operator_8_false_7_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_7_acc_nl);
  assign CONVOLUTION_LOOP_for_for_for_if_2_equal_tmp = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6
      == (operator_8_false_7_acc_tmp[4:0]);
  assign nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6
      + 5'b00001;
  assign CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2[4:0];
  assign nl_operator_8_false_7_acc_tmp = conv_u2s_8_9(n_h_out_lpi_1_dfm) + 9'b111111111;
  assign operator_8_false_7_acc_tmp = nl_operator_8_false_7_acc_tmp[8:0];
  assign nl_operator_8_false_8_acc_nl = ({1'b1 , CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2})
      + 4'b0001;
  assign operator_8_false_8_acc_nl = nl_operator_8_false_8_acc_nl[3:0];
  assign operator_8_false_8_acc_itm_3_1 = readslicef_4_1_3(operator_8_false_8_acc_nl);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2 = CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_4
      + 3'b001;
  assign CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2[2:0];
  assign CONVOLUTION_LOOP_for_for_for_for_not_2310_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0;
  assign CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_4 = MUX_v_3_2_2(3'b000,
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2, CONVOLUTION_LOOP_for_for_for_for_not_2310_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp = CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_4
      == (operator_8_false_4_acc_tmp[2:0]);
  assign exit_CONVOLUTION_LOOP_for_for_for_for_sva_5 = ~((~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp
      & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_cse_sva_1)) | (operator_8_false_4_acc_tmp[8]));
  assign nl_operator_8_false_4_acc_tmp = conv_u2s_8_9(conf_info_crt_sva_231_0[103:96])
      + 9'b111111111;
  assign operator_8_false_4_acc_tmp = nl_operator_8_false_4_acc_tmp[8:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_if_nor_cse_sva_1 = ~((operator_8_false_4_acc_tmp[7:3]!=5'b00000));
  assign nl_operator_8_false_9_acc_nl = ({1'b1 , CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2})
      + 4'b0001;
  assign operator_8_false_9_acc_nl = nl_operator_8_false_9_acc_nl[3:0];
  assign operator_8_false_9_acc_itm_3_1 = readslicef_4_1_3(operator_8_false_9_acc_nl);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2 = CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_5
      + 3'b001;
  assign CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2[2:0];
  assign CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_4_nl
      = lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2 & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0);
  assign CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_5 = MUX_v_3_2_2(3'b000,
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2, CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_4_nl);
  assign or_490_nl = and_769_cse | or_tmp_405;
  assign CONVOLUTION_LOOP_for_mux_1_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0,
      exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1, or_490_nl);
  assign exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4 = CONVOLUTION_LOOP_for_mux_1_nl &
      exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4;
  assign CONVOLUTION_LOOP_for_for_mux_1_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0,
      exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1, or_tmp_405);
  assign exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4 = CONVOLUTION_LOOP_for_for_mux_1_nl
      & exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3;
  assign exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3 = (~(operator_8_false_7_acc_itm_4_1
      & ((~(CONVOLUTION_LOOP_for_for_for_if_2_equal_tmp & (operator_8_false_7_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_7_acc_tmp[8])))) & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1;
  assign exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1 = ~(operator_8_false_9_acc_itm_3_1
      & ((~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_cse_sva_1))
      | (operator_8_false_4_acc_tmp[8])));
  assign CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp = CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_5
      == (operator_8_false_4_acc_tmp[2:0]);
  assign CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_and_1_tmp = lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2
      & lfst_exit_CONVOLUTION_LOOP_for_lpi_2;
  assign nl_BATCH_LOOP_acc_1_tmp = conv_u2u_4_5(BATCH_LOOP_b_4_0_sva_3_0) + 5'b00001;
  assign BATCH_LOOP_acc_1_tmp = nl_BATCH_LOOP_acc_1_tmp[4:0];
  assign BATCH_LOOP_if_2_equal_tmp = BATCH_LOOP_b_4_0_sva_3_0 == (operator_8_false_11_acc_tmp[3:0]);
  assign exit_BATCH_LOOP_sva_2 = ~((~(BATCH_LOOP_if_2_equal_tmp & (operator_8_false_11_acc_tmp[7:4]==4'b0000)))
      | (operator_8_false_11_acc_tmp[8]));
  assign exit_STORE_LOOP_lpi_2_dfm_1 = (~ operator_16_false_1_acc_itm_7_1) | exit_STORE_LOOP_sva_3;
  assign nl_operator_8_false_11_acc_tmp = conv_u2s_8_9(conf_info_crt_sva_231_0[231:224])
      + 9'b111111111;
  assign operator_8_false_11_acc_tmp = nl_operator_8_false_11_acc_tmp[8:0];
  assign nl_operator_16_false_1_acc_nl = conv_u2s_7_8(STORE_LOOP_i_13_0_sva_2[13:7])
      + 8'b10101111;
  assign operator_16_false_1_acc_nl = nl_operator_16_false_1_acc_nl[7:0];
  assign operator_16_false_1_acc_itm_7_1 = readslicef_8_1_7(operator_16_false_1_acc_nl);
  assign nl_STORE_LOOP_i_13_0_sva_2 = STORE_LOOP_i_13_0_lpi_2 + 14'b00000000000001;
  assign STORE_LOOP_i_13_0_sva_2 = nl_STORE_LOOP_i_13_0_sva_2[13:0];
  assign STORE_LOOP_if_equal_tmp = STORE_LOOP_i_13_0_lpi_2 == (operator_16_false_acc_tmp[13:0]);
  assign exit_STORE_LOOP_sva_3 = ~((~(STORE_LOOP_if_equal_tmp & (operator_16_false_acc_tmp[15:14]==2'b00)))
      | (operator_16_false_acc_tmp[16]));
  assign nl_operator_16_false_acc_tmp = conv_u2s_16_17(dma_write_data_length_sva)
      + 17'b11111111111111111;
  assign operator_16_false_acc_tmp = nl_operator_16_false_acc_tmp[16:0];
  assign STORE_LOOP_and_34_ssc_1 = exit_CONVOLUTION_LOOP_lpi_2_dfm_2_1 & STORE_LOOP_equal_tmp_2_1;
  assign STORE_LOOP_equal_tmp_4 = lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0 & lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1
      & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1);
  assign BATCH_LOOP_BATCH_LOOP_or_1_cse_1 = plm_out_data_rsci_bawt | (~(CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3 & lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2
      & (~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1 | lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0))
      & BATCH_LOOP_stage_v_3));
  assign BATCH_LOOP_BATCH_LOOP_or_2_cse_1 = dma_write_chnl_rsci_bawt | (~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_2
      & lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_0 & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_1)
      & BATCH_LOOP_stage_v_4));
  assign CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_mx0 = MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1,
      CONVOLUTION_LOOP_for_for_for_y_lpi_2, and_dcpl_150);
  assign CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_mx0 = MUX_v_8_2_2((z_out_11_16_0[7:0]),
      CONVOLUTION_LOOP_for_for_for_x_lpi_2, and_dcpl_150);
  assign nl_CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6
      * (conf_info_crt_sva_231_0[7:0]);
  assign CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1[7:0];
  assign nl_operator_16_false_acc_nl = conv_u2u_6_7(z_out_12[15:10]) + 7'b1001111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[6:0];
  assign exit_LOAD_LOOP_lpi_2_dfm_1 = (~ (readslicef_7_1_6(operator_16_false_acc_nl)))
      | LOAD_LOOP_LOAD_LOOP_if_and_tmp;
  assign nl_PADDING_LOOP_chan_5_0_sva_2 = conv_u2u_5_6(PADDING_LOOP_chan_5_0_lpi_2_4_0)
      + 6'b000001;
  assign PADDING_LOOP_chan_5_0_sva_2 = nl_PADDING_LOOP_chan_5_0_sva_2[5:0];
  assign or_639_nl = (~ PADDING_LOOP_for_if_equal_tmp) | (operator_8_false_2_acc_tmp[8:5]!=4'b0000)
      | and_dcpl_79;
  assign mux_477_nl = MUX_s_1_2_2(and_dcpl_79, or_639_nl, operator_8_false_2_acc_itm_4_1);
  assign PADDING_LOOP_mux_1_nl = MUX_s_1_2_2(exit_PADDING_LOOP_lpi_2_dfm_mx0w0, exit_PADDING_LOOP_lpi_2_dfm,
      mux_477_nl);
  assign exit_PADDING_LOOP_lpi_2_dfm_3 = PADDING_LOOP_mux_1_nl & exit_PADDING_LOOP_for_lpi_2_dfm_4;
  assign STORE_LOOP_and_tmp_1 = (~ exit_BATCH_LOOP_sva_2) & exit_STORE_LOOP_lpi_2_dfm_1;
  assign STORE_LOOP_equal_tmp_5 = lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1 & lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1
      & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0);
  assign STORE_LOOP_equal_tmp_6 = lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1 & (~(lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0
      | lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1));
  assign STORE_LOOP_or_tmp_2 = (lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0 & lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1
      & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1)) | (lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0
      & lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1 & lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1);
  assign CONVOLUTION_LOOP_for_and_tmp_1 = (~ exit_CONVOLUTION_LOOP_sva_2) & exit_CONVOLUTION_LOOP_for_lpi_2_dfm_4;
  assign PADDING_LOOP_for_and_tmp_1 = (~ exit_PADDING_LOOP_sva_2) & exit_PADDING_LOOP_for_lpi_2_dfm_4;
  assign STORE_LOOP_and_1_m1c_1 = (~ exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1)
      & STORE_LOOP_equal_tmp_2_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_5_tmp_1 = (~ exit_CONVOLUTION_LOOP_for_for_for_for_sva_5)
      & exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1;
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_6_nl = (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0)
      & exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1;
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_7_nl = exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0
      & exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1;
  assign CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_3 = MUX1HOT_v_8_3_2(z_out_13, CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2,
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1, {(~ exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1)
      , CONVOLUTION_LOOP_for_for_for_for_for_and_6_nl , CONVOLUTION_LOOP_for_for_for_for_for_and_7_nl});
  assign nl_CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1 = conv_u2u_2_5(CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[4:3])
      + CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6;
  assign CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1 = nl_CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1[4:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1 = CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6
      + conv_u2u_4_5(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6[4:1]);
  assign CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1 = nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[4:0];
  assign CONVOLUTION_LOOP_for_for_for_asn_3570 = (~(CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3572 = CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3574 = CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3576 = (~(CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3578 = CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3580 = CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3582 = (~(CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3584 = CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3586 = CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3588 = (~(CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3590 = CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3592 = CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3594 = (~(CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3596 = CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3598 = CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3600 = (~(CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3602 = CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3604 = CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3606 = (~(CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3608 = CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3610 = CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3612 = (~(CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3614 = CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3616 = CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3618 = (~(CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3620 = CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3622 = CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3624 = (~(CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3626 = CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3628 = CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3630 = (~(CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3632 = CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3634 = CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3636 = (~(CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3638 = CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3640 = CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3642 = (~(CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3644 = CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3646 = CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3648 = (~(CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3650 = CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3652 = CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3654 = (~(CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3656 = CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3658 = CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3660 = (~(CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3662 = CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3664 = CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3666 = (~(CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3668 = CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3670 = CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3672 = (~(CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3674 = CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3676 = CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3678 = (~(CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3680 = CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3682 = CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3684 = (~(CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3686 = CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3688 = CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3690 = (~(CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3692 = CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3694 = CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3696 = (~(CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3698 = CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3700 = CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3702 = (~(CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3704 = CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3706 = CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3708 = (~(CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3710 = CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3712 = CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3714 = (~(CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3716 = CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3718 = CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3720 = (~(CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3722 = CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3724 = CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3726 = (~(CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3728 = CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3730 = CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3732 = (~(CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3734 = CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3736 = CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3738 = (~(CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3740 = CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3742 = CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3744 = (~(CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3746 = CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3748 = CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3750 = (~(CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3752 = CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3754 = CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3756 = (~(CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3758 = CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3760 = CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3762 = (~(CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3764 = CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3766 = CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3768 = (~(CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3770 = CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3772 = CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3774 = (~(CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3776 = CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3778 = CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3780 = (~(CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3782 = CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3784 = CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3786 = (~(CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3788 = CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3790 = CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3792 = (~(CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3794 = CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3796 = CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3798 = (~(CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3800 = CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3802 = CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3804 = (~(CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3806 = CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3808 = CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3810 = (~(CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3812 = CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3814 = CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3816 = (~(CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3818 = CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3820 = CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3822 = (~(CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3824 = CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3826 = CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3828 = (~(CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3830 = CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3832 = CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3834 = (~(CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3836 = CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3838 = CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3840 = (~(CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3842 = CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3844 = CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3846 = (~(CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3848 = CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3850 = CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3852 = (~(CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3854 = CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3856 = CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3858 = (~(CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3860 = CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3862 = CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3864 = (~(CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3866 = CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3868 = CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3870 = (~(CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3872 = CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3874 = CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3876 = (~(CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3878 = CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3880 = CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3882 = (~(CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3884 = CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3886 = CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3888 = (~(CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3890 = CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3892 = CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3894 = (~(CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3896 = CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3898 = CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3900 = (~(CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3902 = CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3904 = CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3906 = (~(CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3908 = CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3910 = CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3912 = (~(CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3914 = CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3916 = CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3918 = (~(CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3920 = CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3922 = CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3924 = (~(CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3926 = CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3928 = CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3930 = (~(CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3932 = CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3934 = CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3936 = (~(CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3938 = CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3940 = CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3942 = (~(CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3944 = CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3946 = CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3948 = (~(CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3950 = CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3952 = CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3954 = (~(CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3956 = CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3958 = CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3960 = (~(CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3962 = CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3964 = CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3966 = (~(CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3968 = CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3970 = CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3972 = (~(CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3974 = CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3976 = CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3978 = (~(CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3980 = CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3982 = CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3984 = (~(CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3986 = CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3988 = CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3990 = (~(CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3992 = CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3994 = CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3996 = (~(CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3998 = CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4000 = CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4002 = (~(CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4004 = CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4006 = CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4008 = (~(CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4010 = CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4012 = CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4014 = (~(CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4016 = CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4018 = CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4020 = (~(CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4022 = CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4024 = CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4026 = (~(CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4028 = CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4030 = CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4032 = (~(CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4034 = CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4036 = CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4038 = (~(CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4040 = CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4042 = CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4044 = (~(CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4046 = CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4048 = CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4050 = (~(CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4052 = CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4054 = CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4056 = (~(CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4058 = CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4060 = CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4062 = (~(CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4064 = CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4066 = CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4068 = (~(CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4070 = CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4072 = CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4074 = (~(CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4076 = CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4078 = CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4080 = (~(CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4082 = CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4084 = CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4086 = (~(CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4088 = CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4090 = CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4092 = (~(CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4094 = CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4096 = CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4098 = (~(CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4100 = CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4102 = CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4104 = (~(CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4106 = CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4108 = CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4110 = (~(CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4112 = CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4114 = CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4116 = (~(CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4118 = CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4120 = CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4122 = (~(CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4124 = CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4126 = CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4128 = (~(CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4130 = CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4132 = CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4134 = (~(CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4136 = CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4138 = CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4140 = (~(CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4142 = CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4144 = CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4146 = (~(CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4148 = CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4150 = CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4152 = (~(CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4154 = CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4156 = CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4158 = (~(CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4160 = CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4162 = CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4164 = (~(CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4166 = CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4168 = CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4170 = (~(CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4172 = CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4174 = CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4176 = (~(CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4178 = CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4180 = CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4182 = (~(CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4184 = CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4186 = CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4188 = (~(CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4190 = CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4192 = CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4194 = (~(CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4196 = CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4198 = CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4200 = (~(CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4202 = CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4204 = CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4206 = (~(CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4208 = CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4210 = CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4212 = (~(CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4214 = CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4216 = CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4218 = (~(CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4220 = CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4222 = CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4224 = (~(CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4226 = CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4228 = CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4230 = (~(CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4232 = CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4234 = CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4236 = (~(CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4238 = CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4240 = CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4242 = (~(CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4244 = CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4246 = CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4248 = (~(CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4250 = CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4252 = CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4254 = (~(CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4256 = CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4258 = CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4260 = (~(CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4262 = CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4264 = CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4266 = (~(CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4268 = CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4270 = CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4272 = (~(CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4274 = CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4276 = CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4278 = (~(CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4280 = CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4282 = CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4284 = (~(CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4286 = CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4288 = CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4290 = (~(CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4292 = CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4294 = CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4296 = (~(CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4298 = CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4300 = CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4302 = (~(CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4304 = CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4306 = CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4308 = (~(CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4310 = CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4312 = CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4314 = (~(CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4316 = CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4318 = CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4320 = (~(CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4322 = CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4324 = CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4326 = (~(CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4328 = CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4330 = CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4332 = (~(CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4334 = CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4336 = CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4338 = (~(CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4340 = CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4342 = CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4344 = (~(CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4346 = CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4348 = CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4350 = (~(CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4352 = CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4354 = CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4356 = (~(CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4358 = CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4360 = CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4362 = (~(CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4364 = CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4366 = CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4368 = (~(CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4370 = CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4372 = CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4374 = (~(CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4376 = CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4378 = CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4380 = (~(CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4382 = CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4384 = CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4386 = (~(CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4388 = CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4390 = CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4392 = (~(CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4394 = CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4396 = CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4398 = (~(CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4400 = CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4402 = CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4404 = (~(CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4406 = CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4408 = CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4410 = (~(CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4412 = CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4414 = CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4416 = (~(CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4418 = CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4420 = CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4422 = (~(CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4424 = CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4426 = CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4428 = (~(CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4430 = CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4432 = CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4434 = (~(CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4436 = CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4438 = CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4440 = (~(CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4442 = CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4444 = CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4446 = (~(CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4448 = CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4450 = CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4452 = (~(CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4454 = CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4456 = CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4458 = (~(CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4460 = CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4462 = CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4464 = (~(CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4466 = CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4468 = CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4470 = (~(CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4472 = CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4474 = CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4476 = (~(CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4478 = CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4480 = CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4482 = (~(CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4484 = CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4486 = CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4488 = (~(CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4490 = CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4492 = CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4494 = (~(CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4496 = CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4498 = CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4500 = (~(CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4502 = CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4504 = CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4506 = (~(CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4508 = CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4510 = CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4512 = (~(CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4514 = CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4516 = CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4518 = (~(CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4520 = CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4522 = CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4524 = (~(CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4526 = CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4528 = CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4530 = (~(CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4532 = CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4534 = CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4536 = (~(CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4538 = CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4540 = CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4542 = (~(CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4544 = CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4546 = CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4548 = (~(CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4550 = CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4552 = CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4554 = (~(CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4556 = CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4558 = CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4560 = (~(CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4562 = CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4564 = CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4566 = (~(CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4568 = CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4570 = CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4572 = (~(CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4574 = CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4576 = CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4578 = (~(CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4580 = CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4582 = CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4584 = (~(CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4586 = CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4588 = CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4590 = (~(CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4592 = CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4594 = CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4596 = (~(CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4598 = CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4600 = CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4602 = (~(CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4604 = CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4606 = CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4608 = (~(CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4610 = CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4612 = CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4614 = (~(CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4616 = CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4618 = CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4620 = (~(CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4622 = CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4624 = CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4626 = (~(CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4628 = CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4630 = CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4632 = (~(CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4634 = CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4636 = CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4638 = (~(CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4640 = CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4642 = CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4644 = (~(CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4646 = CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4648 = CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4650 = (~(CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4652 = CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4654 = CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4656 = (~(CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4658 = CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4660 = CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4662 = (~(CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4664 = CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4666 = CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4668 = (~(CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4670 = CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4672 = CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4674 = (~(CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4676 = CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4678 = CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4680 = (~(CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4682 = CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4684 = CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4686 = (~(CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4688 = CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4690 = CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4692 = (~(CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4694 = CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4696 = CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4698 = (~(CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4700 = CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4702 = CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4704 = (~(CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4706 = CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4708 = CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4710 = (~(CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4712 = CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4714 = CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4716 = (~(CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4718 = CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4720 = CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4722 = (~(CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4724 = CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4726 = CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4728 = (~(CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4730 = CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4732 = CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4734 = (~(CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4736 = CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4738 = CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4740 = (~(CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4742 = CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4744 = CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4746 = (~(CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4748 = CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4750 = CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4752 = (~(CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4754 = CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4756 = CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4758 = (~(CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4760 = CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4762 = CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4764 = (~(CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4766 = CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4768 = CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4770 = (~(CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4772 = CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4774 = CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4776 = (~(CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4778 = CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4780 = CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4782 = (~(CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4784 = CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4786 = CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4788 = (~(CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4790 = CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4792 = CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4794 = (~(CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4796 = CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4798 = CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4800 = (~(CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4802 = CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4804 = CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4806 = (~(CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4808 = CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4810 = CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4812 = (~(CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4814 = CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4816 = CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4818 = (~(CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4820 = CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4822 = CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4824 = (~(CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4826 = CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4828 = CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4830 = (~(CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4832 = CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4834 = CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4836 = (~(CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4838 = CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4840 = CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4842 = (~(CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4844 = CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4846 = CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4848 = (~(CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4850 = CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4852 = CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4854 = (~(CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4856 = CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4858 = CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4860 = (~(CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4862 = CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4864 = CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4866 = (~(CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4868 = CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4870 = CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4872 = (~(CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4874 = CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4876 = CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4878 = (~(CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4880 = CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4882 = CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4884 = (~(CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4886 = CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4888 = CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4890 = (~(CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4892 = CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4894 = CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4896 = (~(CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4898 = CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4900 = CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4902 = (~(CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4904 = CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4906 = CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4908 = (~(CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4910 = CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4912 = CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4914 = (~(CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4916 = CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4918 = CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4920 = (~(CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4922 = CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4924 = CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4926 = (~(CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4928 = CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4930 = CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4932 = (~(CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4934 = CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4936 = CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4938 = (~(CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4940 = CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4942 = CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4944 = (~(CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4946 = CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4948 = CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4950 = (~(CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4952 = CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4954 = CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4956 = (~(CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4958 = CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4960 = CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4962 = (~(CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4964 = CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4966 = CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4968 = (~(CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4970 = CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4972 = CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4974 = (~(CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4976 = CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4978 = CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4980 = (~(CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4982 = CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4984 = CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4986 = (~(CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4988 = CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4990 = CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4992 = (~(CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4994 = CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4996 = CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4998 = (~(CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5000 = CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5002 = CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5004 = (~(CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5006 = CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5008 = CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5010 = (~(CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5012 = CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5014 = CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5016 = (~(CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5018 = CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5020 = CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5022 = (~(CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5024 = CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5026 = CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5028 = (~(CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5030 = CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5032 = CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5034 = (~(CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5036 = CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5038 = CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5040 = (~(CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5042 = CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5044 = CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5046 = (~(CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5048 = CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5050 = CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5052 = (~(CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5054 = CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5056 = CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5058 = (~(CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5060 = CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5062 = CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5064 = (~(CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5066 = CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5068 = CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5070 = (~(CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5072 = CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5074 = CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5076 = (~(CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5078 = CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5080 = CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5082 = (~(CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5084 = CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5086 = CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5088 = (~(CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5090 = CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5092 = CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5094 = (~(CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5096 = CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5098 = CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5100 = (~(CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5102 = CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5104 = CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5106 = (~(CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5108 = CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5110 = CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5112 = (~(CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5114 = CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5116 = CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5118 = (~(CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5120 = CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5122 = CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5124 = (~(CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5126 = CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5128 = CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5130 = (~(CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5132 = CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5134 = CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5136 = (~(CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5138 = CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5140 = CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5142 = (~(CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5144 = CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5146 = CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5148 = (~(CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5150 = CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5152 = CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5154 = (~(CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5156 = CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5158 = CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5160 = (~(CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5162 = CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5164 = CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5166 = (~(CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5168 = CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5170 = CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5172 = (~(CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5174 = CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5176 = CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5178 = (~(CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5180 = CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5182 = CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5184 = (~(CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5186 = CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5188 = CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5190 = (~(CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5192 = CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5194 = CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5196 = (~(CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5198 = CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5200 = CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5202 = (~(CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5204 = CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5206 = CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5208 = (~(CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5210 = CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5212 = CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5214 = (~(CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5216 = CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5218 = CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5220 = (~(CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5222 = CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5224 = CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5226 = (~(CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5228 = CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5230 = CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5232 = (~(CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5234 = CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5236 = CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5238 = (~(CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5240 = CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5242 = CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5244 = (~(CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5246 = CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5248 = CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5250 = (~(CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5252 = CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5254 = CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5256 = (~(CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5258 = CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5260 = CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5262 = (~(CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5264 = CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5266 = CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5268 = (~(CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5270 = CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5272 = CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5274 = (~(CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5276 = CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5278 = CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5280 = (~(CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5282 = CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5284 = CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5286 = (~(CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5288 = CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5290 = CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5292 = (~(CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5294 = CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5296 = CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5298 = (~(CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5300 = CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5302 = CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5304 = (~(CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5306 = CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5308 = CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5310 = (~(CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5312 = CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5314 = CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5316 = (~(CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5318 = CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5320 = CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5322 = (~(CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5324 = CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5326 = CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5328 = (~(CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5330 = CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5332 = CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5334 = (~(CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5336 = CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5338 = CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5340 = (~(CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5342 = CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5344 = CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5346 = (~(CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5348 = CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5350 = CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5352 = (~(CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5354 = CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5356 = CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5358 = (~(CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5360 = CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5362 = CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5364 = (~(CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5366 = CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5368 = CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5370 = (~(CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5372 = CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5374 = CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5376 = (~(CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5378 = CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5380 = CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5382 = (~(CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5384 = CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5386 = CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5388 = (~(CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5390 = CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5392 = CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5394 = (~(CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5396 = CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5398 = CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5400 = (~(CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5402 = CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5404 = CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5406 = (~(CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5408 = CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5410 = CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5412 = (~(CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5414 = CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5416 = CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5418 = (~(CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5420 = CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5422 = CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5424 = (~(CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5426 = CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5428 = CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5430 = (~(CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5432 = CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5434 = CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5436 = (~(CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5438 = CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5440 = CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5442 = (~(CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5444 = CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5446 = CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5448 = (~(CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5450 = CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5452 = CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5454 = (~(CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5456 = CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5458 = CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5460 = (~(CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5462 = CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5464 = CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5466 = (~(CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5468 = CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5470 = CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5472 = (~(CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5474 = CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5476 = CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5478 = (~(CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5480 = CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5482 = CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5484 = (~(CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5486 = CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5488 = CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5490 = (~(CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5492 = CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5494 = CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5496 = (~(CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5498 = CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5500 = CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5502 = (~(CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5504 = CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5506 = CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5508 = (~(CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5510 = CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5512 = CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign STORE_LOOP_asn_3330 = exit_CONVOLUTION_LOOP_for_for_for_for_for_lpi_2_dfm_1
      & STORE_LOOP_equal_tmp_2_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      = ~((~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[56]) | CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1))
      | CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1);
  assign BATCH_LOOP_and_6_tmp = BATCH_LOOP_stage_v & (~(BATCH_LOOP_stage_v_1 & (~
      BATCH_LOOP_and_4_tmp))) & BATCH_LOOP_stage_0_1 & (plm_f_data_rsci_bawt | (~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1
      & (~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2 | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0))
      & BATCH_LOOP_stage_v_2))) & (plm_in_data_rsci_bawt | (~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1
      & lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0 & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2)
      & BATCH_LOOP_stage_v_2))) & BATCH_LOOP_BATCH_LOOP_or_1_cse_1 & BATCH_LOOP_BATCH_LOOP_or_2_cse_1;
  assign BATCH_LOOP_and_4_tmp = BATCH_LOOP_stage_v_1 & (~(BATCH_LOOP_stage_v_2 &
      or_dcpl_56)) & BATCH_LOOP_stage_0_2 & (dma_read_ctrl_rsci_bawt | (~((reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse
      & (~(reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse)))
      | (~(reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse
      | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse))))) & (dma_read_chnl_rsci_bawt
      | (~(reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse & (~(reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse
      | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse))))) & (dma_read_chnl_rsci_bawt
      | (~(PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1 & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse
      & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse))))
      & (dma_write_ctrl_rsci_bawt | (~(exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1 & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse
      & (~(reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse)))))
      & BATCH_LOOP_BATCH_LOOP_or_1_cse_1 & BATCH_LOOP_BATCH_LOOP_or_2_cse_1;
  assign or_2_cse = (~ BATCH_LOOP_stage_v_4) | dma_write_chnl_rsci_bawt | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_2)
      | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_0) | lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_1;
  assign or_tmp_16 = dma_write_chnl_rsci_bawt | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_2)
      | lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_1 | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_0);
  assign or_tmp_17 = BATCH_LOOP_stage_0 | (~ or_tmp_16);
  assign or_1098_cse = (~ STORE_LOOP_if_equal_tmp) | (operator_16_false_acc_tmp[16:14]!=3'b000);
  assign nand_109_cse = ~(BATCH_LOOP_stage_v_3 & BATCH_LOOP_stage_0_4);
  assign nor_21_cse = ~((operator_16_false_acc_tmp[16:14]!=3'b000) | (~ STORE_LOOP_if_equal_tmp));
  assign or_1096_cse = (operator_8_false_11_acc_tmp[8:4]!=5'b00000) | (~ BATCH_LOOP_if_2_equal_tmp);
  assign and_831_cse = or_1096_cse & BATCH_LOOP_stage_0;
  assign or_131_cse = (~ lfst_exit_STORE_LOOP_lpi_2_1) | lfst_exit_STORE_LOOP_lpi_2_2
      | (~ lfst_exit_STORE_LOOP_lpi_2_0) | exitL_exit_STORE_LOOP_sva;
  assign or_156_cse = lfst_exit_STORE_LOOP_lpi_2_1 | (~ lfst_exit_STORE_LOOP_lpi_2_2)
      | lfst_exit_STORE_LOOP_lpi_2_0 | exitL_exit_STORE_LOOP_sva;
  assign not_tmp_164 = ~(BATCH_LOOP_stage_0_3 & BATCH_LOOP_stage_v_2);
  assign or_tmp_284 = (~ STORE_LOOP_or_2336_tmp) | (~ STORE_LOOP_STORE_LOOP_or_tmp)
      | STORE_LOOP_or_2335_tmp;
  assign nand_90_nl = ~((~(or_1098_cse & BATCH_LOOP_stage_0)) & or_tmp_16);
  assign mux_316_itm = MUX_s_1_2_2((~ or_tmp_16), nand_90_nl, operator_16_false_1_acc_itm_7_1);
  assign mux_560_nl = MUX_s_1_2_2(or_tmp_17, mux_316_itm, or_306_cse);
  assign mux_319_nl = MUX_s_1_2_2(mux_560_nl, or_tmp_17, and_830_cse);
  assign mux_320_nl = MUX_s_1_2_2(mux_319_nl, or_tmp_17, or_tmp_284);
  assign mux_541_nl = MUX_s_1_2_2(or_tmp_17, mux_316_itm, or_306_cse);
  assign mux_318_nl = MUX_s_1_2_2(mux_541_nl, or_tmp_17, or_81_cse);
  assign mux_321_nl = MUX_s_1_2_2(mux_320_nl, mux_318_nl, or_214_cse);
  assign mux_322_nl = MUX_s_1_2_2(or_tmp_17, mux_321_nl, BATCH_LOOP_and_6_tmp);
  assign and_dcpl_16 = ~(mux_322_nl | (~ BATCH_LOOP_stage_v_4) | BATCH_LOOP_stage_0_4
      | BATCH_LOOP_stage_0_3 | BATCH_LOOP_stage_0_1 | BATCH_LOOP_stage_0_2);
  assign or_dcpl_28 = (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2) | lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1
      | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0) | nand_109_cse;
  assign and_dcpl_19 = lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_0 & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_1)
      & lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_2;
  assign and_dcpl_20 = and_dcpl_19 & (~ dma_write_chnl_rsci_bawt) & BATCH_LOOP_stage_v_4;
  assign or_tmp_293 = (~ STORE_LOOP_STORE_LOOP_or_tmp) | STORE_LOOP_or_2336_tmp |
      STORE_LOOP_or_2335_tmp;
  assign or_1104_nl = (~(STORE_LOOP_STORE_LOOP_or_tmp | STORE_LOOP_or_2335_tmp))
      | and_830_cse;
  assign or_334_nl = (~(lfst_exit_STORE_LOOP_lpi_2_2 | lfst_exit_STORE_LOOP_lpi_2_1))
      | exitL_exit_STORE_LOOP_sva;
  assign mux_tmp_319 = MUX_s_1_2_2(or_1104_nl, or_334_nl, or_214_cse);
  assign and_dcpl_22 = BATCH_LOOP_stage_0_3 & BATCH_LOOP_stage_v_2;
  assign and_dcpl_23 = and_dcpl_22 & lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2;
  assign not_tmp_186 = ~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2 | and_dcpl_20);
  assign nor_286_nl = ~(BATCH_LOOP_stage_v_3 | and_dcpl_20);
  assign or_337_nl = (~ BATCH_LOOP_stage_v_3) | lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0
      | plm_out_data_rsci_bawt | (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3)
      | (~ CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3)
      | lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1;
  assign mux_327_nl = MUX_s_1_2_2(not_tmp_186, or_2_cse, or_337_nl);
  assign mux_tmp_321 = MUX_s_1_2_2(nor_286_nl, mux_327_nl, BATCH_LOOP_stage_0_4);
  assign and_dcpl_32 = BATCH_LOOP_stage_v_3 & BATCH_LOOP_stage_0_4;
  assign and_dcpl_33 = lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2 & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1);
  assign and_dcpl_45 = BATCH_LOOP_and_4_tmp & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse);
  assign and_dcpl_48 = BATCH_LOOP_and_4_tmp & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse;
  assign and_dcpl_55 = and_dcpl_22 & (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2);
  assign and_dcpl_65 = and_dcpl_19 & dma_write_chnl_rsci_bawt & BATCH_LOOP_stage_v_4;
  assign or_1078_cse = (~ PADDING_LOOP_for_for_aelse_1_acc_itm_9_1) | (z_out_1_8_0[8])
      | (z_out_3[8]) | (~ (z_out_2[9]));
  assign or_tmp_314 = (or_1078_cse & lfst_exit_STORE_LOOP_lpi_2_0) | lfst_exit_STORE_LOOP_lpi_2_2
      | (~ lfst_exit_STORE_LOOP_lpi_2_1) | exitL_exit_STORE_LOOP_sva;
  assign nand_tmp_29 = (or_1078_cse & STORE_LOOP_or_2336_tmp) | STORE_LOOP_STORE_LOOP_or_tmp
      | (~ STORE_LOOP_or_2335_tmp) | and_830_cse;
  assign and_dcpl_69 = and_dcpl_48 & (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse)
      & ((~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse) | PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1);
  assign and_dcpl_74 = and_dcpl_45 & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse &
      (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse) & exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1;
  assign or_376_nl = (~ lfst_exit_STORE_LOOP_lpi_2_2) | lfst_exit_STORE_LOOP_lpi_2_0
      | lfst_exit_STORE_LOOP_lpi_2_1;
  assign mux_339_nl = MUX_s_1_2_2(or_tmp_293, or_376_nl, BATCH_LOOP_asn_itm_1);
  assign or_375_nl = exit_BATCH_LOOP_lpi_2_dfm_2_1 | BATCH_LOOP_asn_itm_1 | (~ STORE_LOOP_STORE_LOOP_or_tmp)
      | STORE_LOOP_or_2336_tmp | STORE_LOOP_or_2335_tmp;
  assign mux_tmp_333 = MUX_s_1_2_2(mux_339_nl, or_375_nl, exitL_exit_STORE_LOOP_sva);
  assign or_dcpl_48 = ~(BATCH_LOOP_and_4_tmp & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse);
  assign or_dcpl_51 = (~ BATCH_LOOP_and_4_tmp) | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse;
  assign or_tmp_367 = plm_in_data_rsci_bawt | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1)
      | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2;
  assign or_tmp_368 = plm_f_data_rsci_bawt | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1)
      | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2;
  assign and_130_nl = or_tmp_368 & mux_tmp_321;
  assign and_129_nl = or_tmp_367 & mux_tmp_321;
  assign mux_tmp_351 = MUX_s_1_2_2(and_130_nl, and_129_nl, lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0);
  assign or_dcpl_56 = (~ mux_tmp_351) | not_tmp_164;
  assign or_tmp_369 = lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0 | plm_out_data_rsci_bawt
      | (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3) | (~ CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3)
      | lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1;
  assign mux_tmp_352 = MUX_s_1_2_2(not_tmp_186, or_2_cse, or_tmp_369);
  assign or_tmp_372 = (~ exit_BATCH_LOOP_lpi_2_dfm_2_1) | exitL_exit_STORE_LOOP_sva;
  assign or_430_nl = STORE_LOOP_or_2336_tmp | STORE_LOOP_STORE_LOOP_or_tmp | STORE_LOOP_or_2335_tmp;
  assign mux_360_nl = MUX_s_1_2_2(or_tmp_372, and_830_cse, or_430_nl);
  assign mux_tmp_354 = MUX_s_1_2_2(mux_360_nl, exitL_exit_STORE_LOOP_sva, or_214_cse);
  assign not_tmp_219 = ~(operator_16_false_1_acc_itm_7_1 & or_1098_cse);
  assign nand_tmp_39 = ~(or_306_cse & not_tmp_219);
  assign or_441_nl = or_tmp_284 | and_830_cse | nand_tmp_39;
  assign or_438_nl = or_81_cse | nand_tmp_39;
  assign mux_tmp_355 = MUX_s_1_2_2(or_441_nl, or_438_nl, or_214_cse);
  assign or_dcpl_60 = ~(mux_tmp_355 & BATCH_LOOP_and_6_tmp);
  assign nor_tmp_142 = ~((~ STORE_LOOP_or_2336_tmp) | STORE_LOOP_STORE_LOOP_or_tmp
      | (~ STORE_LOOP_or_2335_tmp));
  assign nand_40_nl = ~(nor_tmp_142 & (~ and_830_cse));
  assign mux_tmp_356 = MUX_s_1_2_2(nand_40_nl, or_131_cse, or_214_cse);
  assign or_446_nl = (operator_8_false_1_acc_tmp[8:6]!=3'b000) | (~ PADDING_LOOP_for_for_if_1_equal_tmp)
      | (operator_8_false_1_acc_tmp[5]) | mux_tmp_356;
  assign mux_tmp_357 = MUX_s_1_2_2(mux_tmp_356, or_446_nl, operator_8_false_3_acc_itm_4_1);
  assign or_dcpl_65 = (operator_8_false_1_acc_tmp[5]) | (~ PADDING_LOOP_for_for_if_1_equal_tmp)
      | (operator_8_false_1_acc_tmp[8:6]!=3'b000);
  assign and_dcpl_79 = or_dcpl_65 & operator_8_false_3_acc_itm_4_1;
  assign nand_43_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_240_cse
      | (operator_8_false_4_acc_tmp[8:3]!=6'b000000))));
  assign mux_tmp_361 = MUX_s_1_2_2(and_765_cse, nand_43_nl, operator_8_false_8_acc_itm_3_1);
  assign or_tmp_405 = and_770_cse | mux_tmp_361;
  assign or_tmp_439 = BATCH_LOOP_stage_0_2 | BATCH_LOOP_stage_0 | BATCH_LOOP_stage_0_1
      | BATCH_LOOP_stage_0_3 | BATCH_LOOP_stage_0_4;
  assign or_tmp_440 = or_tmp_439 | (~(BATCH_LOOP_stage_v_4 & or_tmp_16));
  assign or_tmp_444 = and_830_cse | (~ or_tmp_440);
  assign or_tmp_449 = (~ or_tmp_16) | BATCH_LOOP_stage_0_4 | BATCH_LOOP_stage_0_3
      | BATCH_LOOP_stage_0_2 | BATCH_LOOP_stage_0_1 | (~ BATCH_LOOP_stage_v_4);
  assign or_tmp_450 = BATCH_LOOP_stage_0 | or_tmp_449;
  assign or_524_nl = and_831_cse | or_tmp_449;
  assign mux_tmp_372 = MUX_s_1_2_2(or_524_nl, or_tmp_449, BATCH_LOOP_acc_1_tmp[4]);
  assign mux_380_nl = MUX_s_1_2_2(or_tmp_450, mux_tmp_372, nor_21_cse);
  assign mux_381_cse_1 = MUX_s_1_2_2(mux_tmp_372, mux_380_nl, operator_16_false_1_acc_itm_7_1);
  assign nor_294_nl = ~(STORE_LOOP_or_2336_tmp | (~ or_tmp_440));
  assign nor_295_nl = ~(lfst_exit_STORE_LOOP_lpi_2_0 | (~ or_tmp_440));
  assign mux_389_nl = MUX_s_1_2_2(nor_294_nl, nor_295_nl, or_214_cse);
  assign or_dcpl_73 = ~(mux_389_nl & BATCH_LOOP_and_6_tmp);
  assign or_tmp_470 = (~ or_tmp_16) | BATCH_LOOP_stage_0_4 | BATCH_LOOP_stage_0_3
      | BATCH_LOOP_stage_0_1;
  assign or_545_cse = BATCH_LOOP_stage_0_2 | BATCH_LOOP_stage_0 | or_tmp_470;
  assign or_546_nl = and_831_cse | or_tmp_470;
  assign mux_tmp_393 = MUX_s_1_2_2(or_546_nl, or_tmp_470, BATCH_LOOP_acc_1_tmp[4]);
  assign or_tmp_473 = BATCH_LOOP_stage_0 | or_tmp_470;
  assign mux_401_nl = MUX_s_1_2_2(or_tmp_473, mux_tmp_393, nor_21_cse);
  assign mux_tmp_395 = MUX_s_1_2_2(mux_tmp_393, mux_401_nl, operator_16_false_1_acc_itm_7_1);
  assign or_548_cse = BATCH_LOOP_stage_0_2 | mux_tmp_395;
  assign or_tmp_492 = (~ or_tmp_16) | BATCH_LOOP_stage_0_4 | BATCH_LOOP_stage_0_3
      | BATCH_LOOP_stage_0_2 | BATCH_LOOP_stage_0_1 | BATCH_LOOP_stage_0 | (~ BATCH_LOOP_stage_v_4);
  assign nor_277_nl = ~(BATCH_LOOP_if_2_equal_tmp | (~ or_tmp_492));
  assign or_71_nl = (operator_8_false_11_acc_tmp[8:4]!=5'b00000);
  assign mux_425_nl = MUX_s_1_2_2(nor_277_nl, or_tmp_492, or_71_nl);
  assign or_tmp_496 = (BATCH_LOOP_acc_1_tmp[4]) | (~ mux_425_nl);
  assign mux_426_nl = MUX_s_1_2_2(or_tmp_492, (~ or_tmp_496), STORE_LOOP_if_equal_tmp);
  assign or_70_nl = (operator_16_false_acc_tmp[16:14]!=3'b000);
  assign mux_427_nl = MUX_s_1_2_2(mux_426_nl, or_tmp_492, or_70_nl);
  assign mux_tmp_421 = MUX_s_1_2_2((~ or_tmp_496), mux_427_nl, operator_16_false_1_acc_itm_7_1);
  assign or_tmp_509 = (~ or_tmp_16) | BATCH_LOOP_stage_0_4 | BATCH_LOOP_stage_0_3
      | BATCH_LOOP_stage_0_1 | BATCH_LOOP_stage_0;
  assign not_tmp_256 = ~(BATCH_LOOP_stage_0_2 | or_tmp_509);
  assign or_596_nl = (~ CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp) | (operator_8_false_4_acc_tmp[8:3]!=6'b000000)
      | not_tmp_256;
  assign mux_441_nl = MUX_s_1_2_2(not_tmp_256, or_596_nl, operator_8_false_8_acc_itm_3_1);
  assign nand_47_nl = ~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & (~(nor_229_cse
      | (operator_8_false_4_acc_tmp[8:3]!=6'b000000) | not_tmp_256)));
  assign mux_tmp_435 = MUX_s_1_2_2(mux_441_nl, nand_47_nl, operator_8_false_9_acc_itm_3_1);
  assign not_tmp_258 = ~(and_830_cse | mux_tmp_435);
  assign or_619_cse = (~ operator_8_false_9_acc_itm_3_1) | CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp;
  assign or_618_cse = operator_8_false_9_acc_itm_3_1 | operator_8_false_8_acc_itm_3_1;
  assign or_617_cse = (operator_8_false_4_acc_tmp[8:3]!=6'b000000);
  assign nor_272_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp | (~(operator_8_false_8_acc_itm_3_1
      & or_tmp_473)));
  assign mux_452_nl = MUX_s_1_2_2(or_tmp_473, nor_272_nl, or_619_cse);
  assign and_165_nl = or_618_cse & or_tmp_473;
  assign mux_tmp_446 = MUX_s_1_2_2(mux_452_nl, and_165_nl, or_617_cse);
  assign nand_72_nl = ~(or_619_cse & (CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp
      | (~ operator_8_false_8_acc_itm_3_1)));
  assign mux_451_nl = MUX_s_1_2_2(nand_72_nl, or_618_cse, or_617_cse);
  assign mux_tmp_447 = MUX_s_1_2_2(mux_tmp_446, mux_451_nl, BATCH_LOOP_stage_0_2);
  assign mux_tmp_468 = MUX_s_1_2_2(or_324_cse, or_156_cse, or_214_cse);
  assign or_dcpl_85 = mux_tmp_468 | (~ BATCH_LOOP_and_6_tmp);
  assign or_dcpl_87 = not_tmp_164 | BATCH_LOOP_asn_itm_2;
  assign or_dcpl_88 = (~ mux_tmp_351) | or_dcpl_87;
  assign not_tmp_275 = ~((~ or_tmp_16) | BATCH_LOOP_stage_0_4 | BATCH_LOOP_stage_0_3
      | BATCH_LOOP_stage_0_2 | BATCH_LOOP_stage_0_1 | BATCH_LOOP_stage_0 | (~ BATCH_LOOP_stage_v_4));
  assign or_652_nl = (~ CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp) | (operator_8_false_4_acc_tmp[8:3]!=6'b000000)
      | not_tmp_275;
  assign mux_478_nl = MUX_s_1_2_2(not_tmp_275, or_652_nl, operator_8_false_8_acc_itm_3_1);
  assign nand_51_nl = ~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & (~(nor_229_cse
      | (operator_8_false_4_acc_tmp[8:3]!=6'b000000) | not_tmp_275)));
  assign mux_tmp_472 = MUX_s_1_2_2(mux_478_nl, nand_51_nl, operator_8_false_9_acc_itm_3_1);
  assign nor_268_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp | (~(operator_8_false_8_acc_itm_3_1
      & or_tmp_450)));
  assign mux_485_nl = MUX_s_1_2_2(or_tmp_450, nor_268_nl, or_619_cse);
  assign and_170_nl = or_618_cse & or_tmp_450;
  assign mux_486_cse = MUX_s_1_2_2(mux_485_nl, and_170_nl, or_617_cse);
  assign not_tmp_291 = ~(or_tmp_439 | (~ or_tmp_16));
  assign and_dcpl_107 = ~((CONVOLUTION_LOOP_for_k_slc_CONVOLUTION_LOOP_for_k_5_0_4_0_3_itm_1[1:0]!=2'b00));
  assign and_dcpl_109 = ~((CONVOLUTION_LOOP_for_k_slc_CONVOLUTION_LOOP_for_k_5_0_4_0_3_itm_1[4:2]!=3'b000));
  assign or_714_nl = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (~ lfst_exit_STORE_LOOP_lpi_2_2)
      | lfst_exit_STORE_LOOP_lpi_2_1 | exitL_exit_STORE_LOOP_sva | (operator_8_false_4_acc_tmp[8:3]!=6'b000000);
  assign mux_516_nl = MUX_s_1_2_2(or_141_cse, or_714_nl, operator_8_false_9_acc_itm_3_1);
  assign nand_54_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_240_cse
      | (~ lfst_exit_STORE_LOOP_lpi_2_2) | lfst_exit_STORE_LOOP_lpi_2_1 | exitL_exit_STORE_LOOP_sva
      | (operator_8_false_4_acc_tmp[8:3]!=6'b000000))));
  assign mux_tmp_510 = MUX_s_1_2_2(mux_516_nl, nand_54_nl, operator_8_false_8_acc_itm_3_1);
  assign or_tmp_625 = and_830_cse | (operator_8_false_4_acc_tmp[8:3]!=6'b000000);
  assign or_726_nl = (~ STORE_LOOP_STORE_LOOP_or_tmp) | STORE_LOOP_or_2335_tmp |
      and_830_cse;
  assign or_724_nl = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (~ STORE_LOOP_STORE_LOOP_or_tmp)
      | STORE_LOOP_or_2335_tmp | or_tmp_625;
  assign mux_518_nl = MUX_s_1_2_2(or_726_nl, or_724_nl, operator_8_false_9_acc_itm_3_1);
  assign nand_55_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_240_cse
      | (~ STORE_LOOP_STORE_LOOP_or_tmp) | STORE_LOOP_or_2335_tmp | or_tmp_625)));
  assign mux_tmp_512 = MUX_s_1_2_2(mux_518_nl, nand_55_nl, operator_8_false_8_acc_itm_3_1);
  assign or_tmp_645 = ((~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2) & lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2
      & lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2 & lfst_exit_CONVOLUTION_LOOP_for_lpi_2)
      | mux_tmp_468;
  assign and_dcpl_128 = mux_tmp_351 & and_dcpl_22;
  assign not_tmp_312 = ~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1 | (~ or_2_cse));
  assign nand_tmp_57 = ~(or_1096_cse & not_tmp_219);
  assign and_dcpl_138 = (conf_info_rsci_idat_mxwt[7:0]==8'b00000001);
  assign or_dcpl_124 = (~ mux_tmp_351) | not_tmp_164 | BATCH_LOOP_asn_itm_2 | (~
      STORE_LOOP_equal_tmp_2_2);
  assign or_dcpl_127 = (~ mux_tmp_351) | or_dcpl_87 | (~(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2
      & STORE_LOOP_equal_tmp_2_2));
  assign and_dcpl_145 = and_dcpl_109 & and_dcpl_107 & BATCH_LOOP_and_4_tmp;
  assign and_dcpl_150 = CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_and_1_tmp & lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2
      & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2);
  assign or_316_cse = (~((~ CONVOLUTION_LOOP_if_equal_tmp) | (operator_8_false_10_acc_tmp[8:5]!=4'b0000)))
      | (CONVOLUTION_LOOP_acc_tmp[5]);
  assign or_tmp_676 = or_2_cse & and_dcpl_33 & lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0
      & and_dcpl_32 & (fsm_output[2]);
  assign or_tmp_685 = or_dcpl_28 & and_dcpl_65 & (fsm_output[2]);
  assign mux_332_nl = MUX_s_1_2_2(nand_tmp_29, or_tmp_314, BATCH_LOOP_asn_itm_1);
  assign or_tmp_693 = (mux_332_nl | (~ BATCH_LOOP_and_6_tmp)) & and_dcpl_69 & (fsm_output[2]);
  assign or_380_nl = (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | (operator_8_false_4_acc_tmp[8:3]!=6'b000000)
      | mux_tmp_333;
  assign mux_341_nl = MUX_s_1_2_2(mux_tmp_333, or_380_nl, operator_8_false_9_acc_itm_3_1);
  assign nand_34_nl = ~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & (~(nor_240_cse
      | (operator_8_false_4_acc_tmp[8:3]!=6'b000000) | mux_tmp_333)));
  assign mux_342_nl = MUX_s_1_2_2(mux_341_nl, nand_34_nl, operator_8_false_8_acc_itm_3_1);
  assign or_tmp_700 = (~(or_316_cse & or_453_cse & (~(and_769_cse | and_770_cse |
      mux_342_nl)) & BATCH_LOOP_and_6_tmp)) & and_dcpl_74 & (fsm_output[2]);
  assign or_tmp_709 = (~ (fsm_output[2])) | (~ mux_tmp_321) | not_tmp_164 | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2)
      | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1 | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0
      | (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_2) | (~ CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2);
  assign or_tmp_714 = (~ (fsm_output[2])) | or_dcpl_48 | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse
      | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse;
  assign or_tmp_715 = (~ (fsm_output[2])) | or_dcpl_51 | (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse)
      | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse;
  assign or_tmp_717 = (~ (fsm_output[2])) | or_dcpl_48 | reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse
      | (~ reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse);
  assign nor_307_nl = ~(or_tmp_293 | or_tmp_444);
  assign nor_308_nl = ~(or_156_cse | (~ or_tmp_440));
  assign mux_390_nl = MUX_s_1_2_2(nor_307_nl, nor_308_nl, or_214_cse);
  assign or_tmp_760 = mux_390_nl & BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign nor_306_cse = ~((CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0!=5'b00000));
  assign nor_303_cse = ~((CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0!=5'b00000));
  assign or_668_cse = (CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0!=5'b00000);
  assign mux_490_cse = MUX_s_1_2_2(mux_381_cse_1, or_tmp_450, and_830_cse);
  assign mux_484_cse = MUX_s_1_2_2(mux_381_cse_1, or_tmp_450, exitL_exit_STORE_LOOP_sva);
  assign mux_561_nl = MUX_s_1_2_2(mux_486_cse, or_tmp_450, and_830_cse);
  assign mux_492_nl = MUX_s_1_2_2(or_tmp_450, mux_561_nl, or_668_cse);
  assign mux_493_nl = MUX_s_1_2_2(mux_492_nl, mux_490_cse, STORE_LOOP_or_2336_tmp);
  assign mux_494_nl = MUX_s_1_2_2(or_tmp_450, mux_493_nl, nor_93_cse);
  assign or_663_nl = nor_306_cse | exitL_exit_STORE_LOOP_sva;
  assign mux_487_nl = MUX_s_1_2_2(mux_486_cse, or_tmp_450, or_663_nl);
  assign mux_488_nl = MUX_s_1_2_2(mux_487_nl, mux_484_cse, lfst_exit_STORE_LOOP_lpi_2_0);
  assign mux_489_nl = MUX_s_1_2_2(or_tmp_450, mux_488_nl, nor_90_cse);
  assign mux_495_nl = MUX_s_1_2_2(mux_494_nl, mux_489_nl, or_214_cse);
  assign or_tmp_801 = mux_495_nl & BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign mux_558_nl = MUX_s_1_2_2(mux_486_cse, or_tmp_450, and_830_cse);
  assign mux_510_nl = MUX_s_1_2_2(mux_558_nl, or_tmp_450, or_668_cse);
  assign mux_511_nl = MUX_s_1_2_2(mux_510_nl, mux_490_cse, STORE_LOOP_or_2336_tmp);
  assign mux_512_nl = MUX_s_1_2_2(or_tmp_450, mux_511_nl, nor_93_cse);
  assign or_689_nl = (CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0!=5'b00000) | exitL_exit_STORE_LOOP_sva;
  assign mux_505_nl = MUX_s_1_2_2(mux_486_cse, or_tmp_450, or_689_nl);
  assign mux_506_nl = MUX_s_1_2_2(mux_505_nl, mux_484_cse, lfst_exit_STORE_LOOP_lpi_2_0);
  assign mux_507_nl = MUX_s_1_2_2(or_tmp_450, mux_506_nl, nor_90_cse);
  assign mux_513_nl = MUX_s_1_2_2(mux_512_nl, mux_507_nl, or_214_cse);
  assign or_tmp_805 = mux_513_nl & BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign or_tmp_841 = mux_tmp_468 & BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign or_tmp_851 = mux_tmp_351 & and_dcpl_22 & (~ STORE_LOOP_equal_tmp_2_2) &
      (fsm_output[2]);
  assign or_tmp_901 = and_dcpl_138 & (fsm_output[1]);
  assign mux_385_nl = MUX_s_1_2_2(or_tmp_450, mux_381_cse_1, STORE_LOOP_STORE_LOOP_or_tmp);
  assign and_139_nl = STORE_LOOP_STORE_LOOP_or_tmp & or_tmp_450;
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, and_139_nl, STORE_LOOP_or_2335_tmp);
  assign nor_167_nl = ~(and_830_cse | (~ STORE_LOOP_or_2336_tmp));
  assign mux_387_nl = MUX_s_1_2_2(or_tmp_450, mux_386_nl, nor_167_nl);
  assign or_116_nl = (~ lfst_exit_STORE_LOOP_lpi_2_2) | exitL_exit_STORE_LOOP_sva;
  assign mux_382_nl = MUX_s_1_2_2(mux_381_cse_1, or_tmp_450, or_116_nl);
  assign and_138_nl = (lfst_exit_STORE_LOOP_lpi_2_2 | exitL_exit_STORE_LOOP_sva)
      & or_tmp_450;
  assign mux_383_nl = MUX_s_1_2_2(mux_382_nl, and_138_nl, lfst_exit_STORE_LOOP_lpi_2_1);
  assign mux_384_nl = MUX_s_1_2_2(or_tmp_450, mux_383_nl, lfst_exit_STORE_LOOP_lpi_2_0);
  assign mux_388_nl = MUX_s_1_2_2(mux_387_nl, mux_384_nl, or_214_cse);
  assign PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1_mx0c1 = mux_388_nl & BATCH_LOOP_and_6_tmp
      & (fsm_output[2]);
  assign and_151_nl = STORE_LOOP_or_2336_tmp & mux_381_cse_1;
  assign mux_397_nl = MUX_s_1_2_2(and_151_nl, or_tmp_450, and_830_cse);
  assign mux_398_nl = MUX_s_1_2_2(or_tmp_450, mux_397_nl, nor_93_cse);
  assign and_150_nl = exitL_exit_STORE_LOOP_sva & or_tmp_450;
  assign mux_395_nl = MUX_s_1_2_2(and_150_nl, mux_484_cse, lfst_exit_STORE_LOOP_lpi_2_0);
  assign mux_396_nl = MUX_s_1_2_2(or_tmp_450, mux_395_nl, nor_90_cse);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, mux_396_nl, or_214_cse);
  assign exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1_mx0c1 = mux_399_nl & BATCH_LOOP_and_6_tmp
      & (fsm_output[2]);
  assign and_155_nl = lfst_exit_STORE_LOOP_lpi_2_0 & mux_tmp_395;
  assign mux_407_nl = MUX_s_1_2_2(and_155_nl, or_tmp_473, or_141_cse);
  assign and_154_nl = STORE_LOOP_or_2336_tmp & or_548_cse;
  assign mux_404_nl = MUX_s_1_2_2(and_154_nl, or_545_cse, and_830_cse);
  assign mux_405_nl = MUX_s_1_2_2(or_545_cse, mux_404_nl, nor_93_cse);
  assign and_153_nl = lfst_exit_STORE_LOOP_lpi_2_0 & or_548_cse;
  assign mux_403_nl = MUX_s_1_2_2(and_153_nl, or_545_cse, or_141_cse);
  assign mux_406_nl = MUX_s_1_2_2(mux_405_nl, mux_403_nl, BATCH_LOOP_asn_itm_1);
  assign mux_408_nl = MUX_s_1_2_2(mux_407_nl, mux_406_nl, BATCH_LOOP_and_4_tmp);
  assign exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1_mx0c1 = mux_408_nl
      & BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign mux_461_nl = MUX_s_1_2_2(mux_tmp_446, mux_tmp_395, lfst_exit_STORE_LOOP_lpi_2_0);
  assign mux_462_nl = MUX_s_1_2_2(mux_461_nl, or_tmp_473, or_141_cse);
  assign mux_457_nl = MUX_s_1_2_2(mux_tmp_447, or_548_cse, STORE_LOOP_or_2336_tmp);
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, or_545_cse, and_830_cse);
  assign mux_459_nl = MUX_s_1_2_2(or_545_cse, mux_458_nl, nor_93_cse);
  assign mux_455_nl = MUX_s_1_2_2(mux_tmp_447, or_548_cse, lfst_exit_STORE_LOOP_lpi_2_0);
  assign mux_456_nl = MUX_s_1_2_2(mux_455_nl, or_545_cse, or_141_cse);
  assign mux_460_nl = MUX_s_1_2_2(mux_459_nl, mux_456_nl, BATCH_LOOP_asn_itm_1);
  assign mux_463_nl = MUX_s_1_2_2(mux_462_nl, mux_460_nl, BATCH_LOOP_and_4_tmp);
  assign CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1
      = mux_463_nl & BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1_mx0c1 = or_tmp_645 &
      BATCH_LOOP_and_6_tmp & (fsm_output[2]);
  assign BATCH_LOOP_stage_v_2_mx0c0 = (fsm_output[1]) | (mux_tmp_351 & and_dcpl_22
      & (~ BATCH_LOOP_and_4_tmp) & (fsm_output[2]));
  assign and_760_nl = (~(or_tmp_368 & BATCH_LOOP_stage_v_2 & BATCH_LOOP_stage_0_3))
      & mux_tmp_352;
  assign and_761_nl = (~(or_tmp_367 & BATCH_LOOP_stage_v_2 & BATCH_LOOP_stage_0_3))
      & mux_tmp_352;
  assign mux_529_nl = MUX_s_1_2_2(and_760_nl, and_761_nl, lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0);
  assign BATCH_LOOP_stage_v_3_mx0c0 = (fsm_output[1]) | (mux_529_nl & and_dcpl_32
      & (fsm_output[2]));
  assign LOAD_LOOP_i_lpi_2_mx0c1 = (~ BATCH_LOOP_asn_itm_1) & BATCH_LOOP_and_4_tmp
      & (fsm_output[2]);
  assign plm_in_data_rsci_d_d = PADDING_LOOP_for_for_mux_rmff;
  assign plm_in_data_rsci_radr_d = CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff;
  assign plm_in_data_rsci_wadr_d = PADDING_LOOP_for_for_index_in_mux_rmff;
  assign plm_in_data_rsci_we_d_pff = plm_in_data_rsci_we_d_iff;
  assign plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign plm_f_data_rsci_d_d = LOAD_LOOP_data_ac_mux_rmff;
  assign plm_f_data_rsci_radr_d = CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff;
  assign plm_f_data_rsci_wadr_d = LOAD_LOOP_i_mux_rmff;
  assign plm_f_data_rsci_we_d_pff = plm_f_data_rsci_we_d_iff;
  assign plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign plm_out_data_rsci_d_d = {CONVOLUTION_LOOP_for_for_for_if_1_mux_5_rmff ,
      CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff , CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff};
  assign plm_out_data_rsci_radr_d = CONVOLUTION_LOOP_for_for_for_index_out_mux_1_rmff;
  assign plm_out_data_rsci_wadr_d = CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff;
  assign plm_out_data_rsci_we_d_pff = plm_out_data_rsci_we_d_iff;
  assign plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign or_dcpl_135 = STORE_LOOP_or_tmp_2 | STORE_LOOP_or_tmp_mx0w0;
  assign or_dcpl_162 = (or_1066_cse & STORE_LOOP_and_10_cse & exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0)
      | ((~ or_tmp_405) & STORE_LOOP_and_9_m1c);
  assign or_dcpl_163 = ((operator_8_false_8_acc_tmp[8:7]==2'b00) & CONVOLUTION_LOOP_for_for_if_equal_tmp
      & (operator_8_false_8_acc_tmp[6:5]==2'b00) & STORE_LOOP_equal_tmp_2_mx0w0 &
      exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4 & exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0)
      | (or_tmp_405 & STORE_LOOP_and_9_m1c);
  assign or_dcpl_168 = (or_1067_cse & STORE_LOOP_and_12_cse & exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0)
      | ((~ mux_tmp_361) & STORE_LOOP_and_11_m1c);
  assign or_dcpl_169 = (CONVOLUTION_LOOP_for_for_for_if_2_equal_tmp & (operator_8_false_7_acc_tmp[8:5]==4'b0000)
      & STORE_LOOP_equal_tmp_2_mx0w0 & exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3
      & exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0) | (mux_tmp_361 & STORE_LOOP_and_11_m1c);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | and_dcpl_20 | or_dcpl_28)) ) begin
      dma_write_chnl_rsci_idat_31_0 <= plm_out_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_rsci_idat_15_0 <= 16'b0000000000000000;
      dma_write_ctrl_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( BATCH_LOOP_and_cse ) begin
      dma_write_ctrl_rsci_idat_15_0 <= z_out;
      dma_write_ctrl_rsci_idat_47_32 <= dma_write_data_length_sva;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_idat_15_0 <= 16'b0000000000000000;
      dma_read_ctrl_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( LOAD_CTRL_LOOP_and_cse ) begin
      dma_read_ctrl_rsci_idat_15_0 <= MUX_v_16_2_2(dma_read_info_index_15_0_lpi_2,
          z_out_6, mux_526_nl);
      dma_read_ctrl_rsci_idat_47_32 <= dma_read_data_length_sva;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
      reg_plm_out_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= 1'b0;
      reg_plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
      reg_plm_f_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= 1'b0;
      reg_plm_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= 1'b0;
      reg_acc_done_rsci_ivld_core_psct_cse <= 1'b0;
      reg_dma_read_ctrl_rsci_ivld_core_psct_cse <= 1'b0;
      reg_conf_info_rsci_irdy_core_psct_cse <= 1'b0;
      plm_out_data_rsci_wadr_d_reg <= 14'b00000000000000;
      plm_out_data_rsci_radr_d_reg <= 14'b00000000000000;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5 <=
          1'b0;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4 <=
          30'b000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3 <=
          1'b0;
      plm_f_data_rsci_wadr_d_reg <= 16'b0000000000000000;
      plm_f_data_rsci_radr_d_reg <= 16'b0000000000000000;
      plm_f_data_rsci_d_d_reg <= 32'b00000000000000000000000000000000;
      plm_in_data_rsci_wadr_d_reg <= 14'b00000000000000;
      plm_in_data_rsci_radr_d_reg <= 14'b00000000000000;
      plm_in_data_rsci_d_d_reg <= 32'b00000000000000000000000000000000;
      BATCH_LOOP_stage_v <= 1'b0;
      BATCH_LOOP_stage_v_4 <= 1'b0;
      BATCH_LOOP_stage_0 <= 1'b0;
      BATCH_LOOP_b_4_0_sva_3_0 <= 4'b0000;
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0 <= 5'b00000;
      exitL_exit_STORE_LOOP_sva <= 1'b0;
      BATCH_LOOP_stage_v_1 <= 1'b0;
      BATCH_LOOP_stage_0_1 <= 1'b0;
      BATCH_LOOP_stage_0_2 <= 1'b0;
      BATCH_LOOP_stage_0_4 <= 1'b0;
      buf_acc_data_17_17_0_sva <= 1'b0;
      buf_acc_data_17_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_0_0_sva <= 1'b0;
      buf_acc_data_0_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_16_0_sva <= 1'b0;
      buf_acc_data_17_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_1_0_sva <= 1'b0;
      buf_acc_data_0_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_15_0_sva <= 1'b0;
      buf_acc_data_17_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_2_0_sva <= 1'b0;
      buf_acc_data_0_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_14_0_sva <= 1'b0;
      buf_acc_data_17_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_3_0_sva <= 1'b0;
      buf_acc_data_0_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_13_0_sva <= 1'b0;
      buf_acc_data_17_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_4_0_sva <= 1'b0;
      buf_acc_data_0_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_12_0_sva <= 1'b0;
      buf_acc_data_17_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_5_0_sva <= 1'b0;
      buf_acc_data_0_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_11_0_sva <= 1'b0;
      buf_acc_data_17_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_6_0_sva <= 1'b0;
      buf_acc_data_0_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_10_0_sva <= 1'b0;
      buf_acc_data_17_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_7_0_sva <= 1'b0;
      buf_acc_data_0_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_9_0_sva <= 1'b0;
      buf_acc_data_17_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_8_0_sva <= 1'b0;
      buf_acc_data_0_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_8_0_sva <= 1'b0;
      buf_acc_data_17_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_9_0_sva <= 1'b0;
      buf_acc_data_0_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_7_0_sva <= 1'b0;
      buf_acc_data_17_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_10_0_sva <= 1'b0;
      buf_acc_data_0_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_6_0_sva <= 1'b0;
      buf_acc_data_17_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_11_0_sva <= 1'b0;
      buf_acc_data_0_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_5_0_sva <= 1'b0;
      buf_acc_data_17_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_12_0_sva <= 1'b0;
      buf_acc_data_0_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_4_0_sva <= 1'b0;
      buf_acc_data_17_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_13_0_sva <= 1'b0;
      buf_acc_data_0_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_3_0_sva <= 1'b0;
      buf_acc_data_17_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_14_0_sva <= 1'b0;
      buf_acc_data_0_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_2_0_sva <= 1'b0;
      buf_acc_data_17_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_15_0_sva <= 1'b0;
      buf_acc_data_0_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_1_0_sva <= 1'b0;
      buf_acc_data_17_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_16_0_sva <= 1'b0;
      buf_acc_data_0_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_17_0_0_sva <= 1'b0;
      buf_acc_data_17_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_17_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_0_17_0_sva <= 1'b0;
      buf_acc_data_0_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_0_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_17_0_sva <= 1'b0;
      buf_acc_data_16_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_0_0_sva <= 1'b0;
      buf_acc_data_1_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_16_0_sva <= 1'b0;
      buf_acc_data_16_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_1_0_sva <= 1'b0;
      buf_acc_data_1_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_15_0_sva <= 1'b0;
      buf_acc_data_16_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_2_0_sva <= 1'b0;
      buf_acc_data_1_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_14_0_sva <= 1'b0;
      buf_acc_data_16_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_3_0_sva <= 1'b0;
      buf_acc_data_1_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_13_0_sva <= 1'b0;
      buf_acc_data_16_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_4_0_sva <= 1'b0;
      buf_acc_data_1_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_12_0_sva <= 1'b0;
      buf_acc_data_16_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_5_0_sva <= 1'b0;
      buf_acc_data_1_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_11_0_sva <= 1'b0;
      buf_acc_data_16_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_6_0_sva <= 1'b0;
      buf_acc_data_1_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_10_0_sva <= 1'b0;
      buf_acc_data_16_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_7_0_sva <= 1'b0;
      buf_acc_data_1_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_9_0_sva <= 1'b0;
      buf_acc_data_16_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_8_0_sva <= 1'b0;
      buf_acc_data_1_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_8_0_sva <= 1'b0;
      buf_acc_data_16_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_9_0_sva <= 1'b0;
      buf_acc_data_1_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_7_0_sva <= 1'b0;
      buf_acc_data_16_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_10_0_sva <= 1'b0;
      buf_acc_data_1_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_6_0_sva <= 1'b0;
      buf_acc_data_16_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_11_0_sva <= 1'b0;
      buf_acc_data_1_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_5_0_sva <= 1'b0;
      buf_acc_data_16_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_12_0_sva <= 1'b0;
      buf_acc_data_1_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_4_0_sva <= 1'b0;
      buf_acc_data_16_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_13_0_sva <= 1'b0;
      buf_acc_data_1_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_3_0_sva <= 1'b0;
      buf_acc_data_16_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_14_0_sva <= 1'b0;
      buf_acc_data_1_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_2_0_sva <= 1'b0;
      buf_acc_data_16_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_15_0_sva <= 1'b0;
      buf_acc_data_1_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_1_0_sva <= 1'b0;
      buf_acc_data_16_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_16_0_sva <= 1'b0;
      buf_acc_data_1_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_16_0_0_sva <= 1'b0;
      buf_acc_data_16_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_16_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_1_17_0_sva <= 1'b0;
      buf_acc_data_1_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_1_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_17_0_sva <= 1'b0;
      buf_acc_data_15_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_0_0_sva <= 1'b0;
      buf_acc_data_2_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_16_0_sva <= 1'b0;
      buf_acc_data_15_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_1_0_sva <= 1'b0;
      buf_acc_data_2_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_15_0_sva <= 1'b0;
      buf_acc_data_15_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_2_0_sva <= 1'b0;
      buf_acc_data_2_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_14_0_sva <= 1'b0;
      buf_acc_data_15_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_3_0_sva <= 1'b0;
      buf_acc_data_2_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_13_0_sva <= 1'b0;
      buf_acc_data_15_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_4_0_sva <= 1'b0;
      buf_acc_data_2_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_12_0_sva <= 1'b0;
      buf_acc_data_15_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_5_0_sva <= 1'b0;
      buf_acc_data_2_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_11_0_sva <= 1'b0;
      buf_acc_data_15_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_6_0_sva <= 1'b0;
      buf_acc_data_2_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_10_0_sva <= 1'b0;
      buf_acc_data_15_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_7_0_sva <= 1'b0;
      buf_acc_data_2_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_9_0_sva <= 1'b0;
      buf_acc_data_15_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_8_0_sva <= 1'b0;
      buf_acc_data_2_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_8_0_sva <= 1'b0;
      buf_acc_data_15_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_9_0_sva <= 1'b0;
      buf_acc_data_2_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_7_0_sva <= 1'b0;
      buf_acc_data_15_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_10_0_sva <= 1'b0;
      buf_acc_data_2_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_6_0_sva <= 1'b0;
      buf_acc_data_15_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_11_0_sva <= 1'b0;
      buf_acc_data_2_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_5_0_sva <= 1'b0;
      buf_acc_data_15_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_12_0_sva <= 1'b0;
      buf_acc_data_2_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_4_0_sva <= 1'b0;
      buf_acc_data_15_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_13_0_sva <= 1'b0;
      buf_acc_data_2_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_3_0_sva <= 1'b0;
      buf_acc_data_15_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_14_0_sva <= 1'b0;
      buf_acc_data_2_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_2_0_sva <= 1'b0;
      buf_acc_data_15_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_15_0_sva <= 1'b0;
      buf_acc_data_2_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_1_0_sva <= 1'b0;
      buf_acc_data_15_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_16_0_sva <= 1'b0;
      buf_acc_data_2_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_15_0_0_sva <= 1'b0;
      buf_acc_data_15_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_15_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_2_17_0_sva <= 1'b0;
      buf_acc_data_2_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_2_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_17_0_sva <= 1'b0;
      buf_acc_data_14_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_0_0_sva <= 1'b0;
      buf_acc_data_3_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_16_0_sva <= 1'b0;
      buf_acc_data_14_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_1_0_sva <= 1'b0;
      buf_acc_data_3_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_15_0_sva <= 1'b0;
      buf_acc_data_14_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_2_0_sva <= 1'b0;
      buf_acc_data_3_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_14_0_sva <= 1'b0;
      buf_acc_data_14_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_3_0_sva <= 1'b0;
      buf_acc_data_3_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_13_0_sva <= 1'b0;
      buf_acc_data_14_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_4_0_sva <= 1'b0;
      buf_acc_data_3_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_12_0_sva <= 1'b0;
      buf_acc_data_14_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_5_0_sva <= 1'b0;
      buf_acc_data_3_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_11_0_sva <= 1'b0;
      buf_acc_data_14_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_6_0_sva <= 1'b0;
      buf_acc_data_3_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_10_0_sva <= 1'b0;
      buf_acc_data_14_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_7_0_sva <= 1'b0;
      buf_acc_data_3_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_9_0_sva <= 1'b0;
      buf_acc_data_14_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_8_0_sva <= 1'b0;
      buf_acc_data_3_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_8_0_sva <= 1'b0;
      buf_acc_data_14_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_9_0_sva <= 1'b0;
      buf_acc_data_3_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_7_0_sva <= 1'b0;
      buf_acc_data_14_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_10_0_sva <= 1'b0;
      buf_acc_data_3_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_6_0_sva <= 1'b0;
      buf_acc_data_14_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_11_0_sva <= 1'b0;
      buf_acc_data_3_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_5_0_sva <= 1'b0;
      buf_acc_data_14_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_12_0_sva <= 1'b0;
      buf_acc_data_3_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_4_0_sva <= 1'b0;
      buf_acc_data_14_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_13_0_sva <= 1'b0;
      buf_acc_data_3_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_3_0_sva <= 1'b0;
      buf_acc_data_14_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_14_0_sva <= 1'b0;
      buf_acc_data_3_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_2_0_sva <= 1'b0;
      buf_acc_data_14_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_15_0_sva <= 1'b0;
      buf_acc_data_3_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_1_0_sva <= 1'b0;
      buf_acc_data_14_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_16_0_sva <= 1'b0;
      buf_acc_data_3_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_14_0_0_sva <= 1'b0;
      buf_acc_data_14_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_14_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_3_17_0_sva <= 1'b0;
      buf_acc_data_3_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_3_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_17_0_sva <= 1'b0;
      buf_acc_data_13_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_0_0_sva <= 1'b0;
      buf_acc_data_4_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_16_0_sva <= 1'b0;
      buf_acc_data_13_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_1_0_sva <= 1'b0;
      buf_acc_data_4_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_15_0_sva <= 1'b0;
      buf_acc_data_13_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_2_0_sva <= 1'b0;
      buf_acc_data_4_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_14_0_sva <= 1'b0;
      buf_acc_data_13_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_3_0_sva <= 1'b0;
      buf_acc_data_4_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_13_0_sva <= 1'b0;
      buf_acc_data_13_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_4_0_sva <= 1'b0;
      buf_acc_data_4_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_12_0_sva <= 1'b0;
      buf_acc_data_13_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_5_0_sva <= 1'b0;
      buf_acc_data_4_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_11_0_sva <= 1'b0;
      buf_acc_data_13_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_6_0_sva <= 1'b0;
      buf_acc_data_4_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_10_0_sva <= 1'b0;
      buf_acc_data_13_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_7_0_sva <= 1'b0;
      buf_acc_data_4_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_9_0_sva <= 1'b0;
      buf_acc_data_13_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_8_0_sva <= 1'b0;
      buf_acc_data_4_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_8_0_sva <= 1'b0;
      buf_acc_data_13_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_9_0_sva <= 1'b0;
      buf_acc_data_4_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_7_0_sva <= 1'b0;
      buf_acc_data_13_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_10_0_sva <= 1'b0;
      buf_acc_data_4_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_6_0_sva <= 1'b0;
      buf_acc_data_13_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_11_0_sva <= 1'b0;
      buf_acc_data_4_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_5_0_sva <= 1'b0;
      buf_acc_data_13_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_12_0_sva <= 1'b0;
      buf_acc_data_4_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_4_0_sva <= 1'b0;
      buf_acc_data_13_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_13_0_sva <= 1'b0;
      buf_acc_data_4_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_3_0_sva <= 1'b0;
      buf_acc_data_13_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_14_0_sva <= 1'b0;
      buf_acc_data_4_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_2_0_sva <= 1'b0;
      buf_acc_data_13_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_15_0_sva <= 1'b0;
      buf_acc_data_4_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_1_0_sva <= 1'b0;
      buf_acc_data_13_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_16_0_sva <= 1'b0;
      buf_acc_data_4_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_13_0_0_sva <= 1'b0;
      buf_acc_data_13_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_13_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_4_17_0_sva <= 1'b0;
      buf_acc_data_4_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_4_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_17_0_sva <= 1'b0;
      buf_acc_data_12_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_0_0_sva <= 1'b0;
      buf_acc_data_5_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_16_0_sva <= 1'b0;
      buf_acc_data_12_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_1_0_sva <= 1'b0;
      buf_acc_data_5_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_15_0_sva <= 1'b0;
      buf_acc_data_12_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_2_0_sva <= 1'b0;
      buf_acc_data_5_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_14_0_sva <= 1'b0;
      buf_acc_data_12_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_3_0_sva <= 1'b0;
      buf_acc_data_5_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_13_0_sva <= 1'b0;
      buf_acc_data_12_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_4_0_sva <= 1'b0;
      buf_acc_data_5_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_12_0_sva <= 1'b0;
      buf_acc_data_12_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_5_0_sva <= 1'b0;
      buf_acc_data_5_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_11_0_sva <= 1'b0;
      buf_acc_data_12_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_6_0_sva <= 1'b0;
      buf_acc_data_5_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_10_0_sva <= 1'b0;
      buf_acc_data_12_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_7_0_sva <= 1'b0;
      buf_acc_data_5_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_9_0_sva <= 1'b0;
      buf_acc_data_12_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_8_0_sva <= 1'b0;
      buf_acc_data_5_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_8_0_sva <= 1'b0;
      buf_acc_data_12_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_9_0_sva <= 1'b0;
      buf_acc_data_5_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_7_0_sva <= 1'b0;
      buf_acc_data_12_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_10_0_sva <= 1'b0;
      buf_acc_data_5_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_6_0_sva <= 1'b0;
      buf_acc_data_12_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_11_0_sva <= 1'b0;
      buf_acc_data_5_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_5_0_sva <= 1'b0;
      buf_acc_data_12_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_12_0_sva <= 1'b0;
      buf_acc_data_5_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_4_0_sva <= 1'b0;
      buf_acc_data_12_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_13_0_sva <= 1'b0;
      buf_acc_data_5_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_3_0_sva <= 1'b0;
      buf_acc_data_12_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_14_0_sva <= 1'b0;
      buf_acc_data_5_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_2_0_sva <= 1'b0;
      buf_acc_data_12_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_15_0_sva <= 1'b0;
      buf_acc_data_5_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_1_0_sva <= 1'b0;
      buf_acc_data_12_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_16_0_sva <= 1'b0;
      buf_acc_data_5_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_12_0_0_sva <= 1'b0;
      buf_acc_data_12_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_12_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_5_17_0_sva <= 1'b0;
      buf_acc_data_5_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_5_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_17_0_sva <= 1'b0;
      buf_acc_data_11_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_0_0_sva <= 1'b0;
      buf_acc_data_6_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_16_0_sva <= 1'b0;
      buf_acc_data_11_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_1_0_sva <= 1'b0;
      buf_acc_data_6_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_15_0_sva <= 1'b0;
      buf_acc_data_11_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_2_0_sva <= 1'b0;
      buf_acc_data_6_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_14_0_sva <= 1'b0;
      buf_acc_data_11_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_3_0_sva <= 1'b0;
      buf_acc_data_6_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_13_0_sva <= 1'b0;
      buf_acc_data_11_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_4_0_sva <= 1'b0;
      buf_acc_data_6_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_12_0_sva <= 1'b0;
      buf_acc_data_11_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_5_0_sva <= 1'b0;
      buf_acc_data_6_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_11_0_sva <= 1'b0;
      buf_acc_data_11_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_6_0_sva <= 1'b0;
      buf_acc_data_6_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_10_0_sva <= 1'b0;
      buf_acc_data_11_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_7_0_sva <= 1'b0;
      buf_acc_data_6_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_9_0_sva <= 1'b0;
      buf_acc_data_11_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_8_0_sva <= 1'b0;
      buf_acc_data_6_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_8_0_sva <= 1'b0;
      buf_acc_data_11_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_9_0_sva <= 1'b0;
      buf_acc_data_6_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_7_0_sva <= 1'b0;
      buf_acc_data_11_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_10_0_sva <= 1'b0;
      buf_acc_data_6_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_6_0_sva <= 1'b0;
      buf_acc_data_11_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_11_0_sva <= 1'b0;
      buf_acc_data_6_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_5_0_sva <= 1'b0;
      buf_acc_data_11_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_12_0_sva <= 1'b0;
      buf_acc_data_6_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_4_0_sva <= 1'b0;
      buf_acc_data_11_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_13_0_sva <= 1'b0;
      buf_acc_data_6_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_3_0_sva <= 1'b0;
      buf_acc_data_11_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_14_0_sva <= 1'b0;
      buf_acc_data_6_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_2_0_sva <= 1'b0;
      buf_acc_data_11_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_15_0_sva <= 1'b0;
      buf_acc_data_6_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_1_0_sva <= 1'b0;
      buf_acc_data_11_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_16_0_sva <= 1'b0;
      buf_acc_data_6_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_11_0_0_sva <= 1'b0;
      buf_acc_data_11_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_11_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_6_17_0_sva <= 1'b0;
      buf_acc_data_6_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_6_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_17_0_sva <= 1'b0;
      buf_acc_data_10_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_0_0_sva <= 1'b0;
      buf_acc_data_7_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_16_0_sva <= 1'b0;
      buf_acc_data_10_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_1_0_sva <= 1'b0;
      buf_acc_data_7_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_15_0_sva <= 1'b0;
      buf_acc_data_10_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_2_0_sva <= 1'b0;
      buf_acc_data_7_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_14_0_sva <= 1'b0;
      buf_acc_data_10_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_3_0_sva <= 1'b0;
      buf_acc_data_7_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_13_0_sva <= 1'b0;
      buf_acc_data_10_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_4_0_sva <= 1'b0;
      buf_acc_data_7_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_12_0_sva <= 1'b0;
      buf_acc_data_10_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_5_0_sva <= 1'b0;
      buf_acc_data_7_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_11_0_sva <= 1'b0;
      buf_acc_data_10_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_6_0_sva <= 1'b0;
      buf_acc_data_7_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_10_0_sva <= 1'b0;
      buf_acc_data_10_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_7_0_sva <= 1'b0;
      buf_acc_data_7_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_9_0_sva <= 1'b0;
      buf_acc_data_10_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_8_0_sva <= 1'b0;
      buf_acc_data_7_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_8_0_sva <= 1'b0;
      buf_acc_data_10_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_9_0_sva <= 1'b0;
      buf_acc_data_7_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_7_0_sva <= 1'b0;
      buf_acc_data_10_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_10_0_sva <= 1'b0;
      buf_acc_data_7_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_6_0_sva <= 1'b0;
      buf_acc_data_10_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_11_0_sva <= 1'b0;
      buf_acc_data_7_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_5_0_sva <= 1'b0;
      buf_acc_data_10_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_12_0_sva <= 1'b0;
      buf_acc_data_7_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_4_0_sva <= 1'b0;
      buf_acc_data_10_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_13_0_sva <= 1'b0;
      buf_acc_data_7_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_3_0_sva <= 1'b0;
      buf_acc_data_10_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_14_0_sva <= 1'b0;
      buf_acc_data_7_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_2_0_sva <= 1'b0;
      buf_acc_data_10_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_15_0_sva <= 1'b0;
      buf_acc_data_7_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_1_0_sva <= 1'b0;
      buf_acc_data_10_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_16_0_sva <= 1'b0;
      buf_acc_data_7_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_10_0_0_sva <= 1'b0;
      buf_acc_data_10_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_10_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_7_17_0_sva <= 1'b0;
      buf_acc_data_7_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_7_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_17_0_sva <= 1'b0;
      buf_acc_data_9_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_17_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_0_0_sva <= 1'b0;
      buf_acc_data_8_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_16_0_sva <= 1'b0;
      buf_acc_data_9_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_1_0_sva <= 1'b0;
      buf_acc_data_8_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_15_0_sva <= 1'b0;
      buf_acc_data_9_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_2_0_sva <= 1'b0;
      buf_acc_data_8_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_14_0_sva <= 1'b0;
      buf_acc_data_9_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_3_0_sva <= 1'b0;
      buf_acc_data_8_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_13_0_sva <= 1'b0;
      buf_acc_data_9_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_4_0_sva <= 1'b0;
      buf_acc_data_8_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_12_0_sva <= 1'b0;
      buf_acc_data_9_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_5_0_sva <= 1'b0;
      buf_acc_data_8_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_11_0_sva <= 1'b0;
      buf_acc_data_9_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_6_0_sva <= 1'b0;
      buf_acc_data_8_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_10_0_sva <= 1'b0;
      buf_acc_data_9_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_7_0_sva <= 1'b0;
      buf_acc_data_8_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_9_0_sva <= 1'b0;
      buf_acc_data_9_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_8_0_sva <= 1'b0;
      buf_acc_data_8_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_8_0_sva <= 1'b0;
      buf_acc_data_9_8_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_8_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_9_0_sva <= 1'b0;
      buf_acc_data_8_9_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_9_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_7_0_sva <= 1'b0;
      buf_acc_data_9_7_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_7_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_10_0_sva <= 1'b0;
      buf_acc_data_8_10_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_10_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_6_0_sva <= 1'b0;
      buf_acc_data_9_6_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_6_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_11_0_sva <= 1'b0;
      buf_acc_data_8_11_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_11_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_5_0_sva <= 1'b0;
      buf_acc_data_9_5_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_5_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_12_0_sva <= 1'b0;
      buf_acc_data_8_12_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_12_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_4_0_sva <= 1'b0;
      buf_acc_data_9_4_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_4_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_13_0_sva <= 1'b0;
      buf_acc_data_8_13_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_13_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_3_0_sva <= 1'b0;
      buf_acc_data_9_3_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_3_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_14_0_sva <= 1'b0;
      buf_acc_data_8_14_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_14_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_2_0_sva <= 1'b0;
      buf_acc_data_9_2_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_2_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_15_0_sva <= 1'b0;
      buf_acc_data_8_15_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_15_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_1_0_sva <= 1'b0;
      buf_acc_data_9_1_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_1_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_16_0_sva <= 1'b0;
      buf_acc_data_8_16_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_16_56_46_sva <= 11'b00000000000;
      buf_acc_data_9_0_0_sva <= 1'b0;
      buf_acc_data_9_0_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_9_0_56_46_sva <= 11'b00000000000;
      buf_acc_data_8_17_0_sva <= 1'b0;
      buf_acc_data_8_17_45_1_sva <= 45'b000000000000000000000000000000000000000000000;
      buf_acc_data_8_17_56_46_sva <= 11'b00000000000;
      CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= and_245_rmff;
      reg_plm_out_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= and_247_rmff;
      reg_plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= and_253_rmff;
      reg_plm_f_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= and_255_rmff;
      reg_plm_in_data_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= and_261_rmff;
      reg_acc_done_rsci_ivld_core_psct_cse <= and_dcpl_16 & (fsm_output[2]);
      reg_dma_read_ctrl_rsci_ivld_core_psct_cse <= mux_tmp_319 & BATCH_LOOP_and_6_tmp
          & (fsm_output[2]);
      reg_conf_info_rsci_irdy_core_psct_cse <= ~((fsm_output[2:1]!=2'b00));
      plm_out_data_rsci_wadr_d_reg <= CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff;
      plm_out_data_rsci_radr_d_reg <= CONVOLUTION_LOOP_for_for_for_index_out_mux_1_rmff;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5 <=
          CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4 <=
          CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3 <=
          CONVOLUTION_LOOP_for_for_for_if_1_mux_5_rmff;
      plm_f_data_rsci_wadr_d_reg <= LOAD_LOOP_i_mux_rmff;
      plm_f_data_rsci_radr_d_reg <= CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff;
      plm_f_data_rsci_d_d_reg <= LOAD_LOOP_data_ac_mux_rmff;
      plm_in_data_rsci_wadr_d_reg <= PADDING_LOOP_for_for_index_in_mux_rmff;
      plm_in_data_rsci_radr_d_reg <= CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff;
      plm_in_data_rsci_d_d_reg <= PADDING_LOOP_for_for_mux_rmff;
      BATCH_LOOP_stage_v <= ~((~(BATCH_LOOP_stage_v & (~((~(mux_tmp_355 & BATCH_LOOP_stage_0))
          & BATCH_LOOP_and_6_tmp)))) & (~(mux_528_nl & BATCH_LOOP_stage_0)) & (fsm_output[2]));
      BATCH_LOOP_stage_v_4 <= ((BATCH_LOOP_stage_v_4 & (~ mux_534_nl)) | (mux_tmp_352
          & and_dcpl_32)) & (fsm_output[2]);
      BATCH_LOOP_stage_0 <= ~((~(BATCH_LOOP_stage_0 & (mux_tmp_355 | (~ BATCH_LOOP_and_6_tmp))))
          & (fsm_output[2]));
      BATCH_LOOP_b_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, STORE_LOOP_mux_37_nl, (fsm_output[2]));
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0 <= MUX_v_5_2_2(CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0,
          CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1, fsm_output[2]);
      exitL_exit_STORE_LOOP_sva <= exitL_exit_STORE_LOOP_sva_mx1 | (~ (fsm_output[2]));
      BATCH_LOOP_stage_v_1 <= ((BATCH_LOOP_stage_v_1 & (~ BATCH_LOOP_and_4_tmp))
          | BATCH_LOOP_and_6_tmp) & (fsm_output[2]);
      BATCH_LOOP_stage_0_1 <= ~((~(PADDING_LOOP_for_for_aelse_mux_nl & (~((~ mux_tmp_355)
          & BATCH_LOOP_and_6_tmp)))) & (fsm_output[2]));
      BATCH_LOOP_stage_0_2 <= BATCH_LOOP_mux_5_nl & (fsm_output[2]);
      BATCH_LOOP_stage_0_4 <= BATCH_LOOP_mux_6_nl & (fsm_output[2]);
      buf_acc_data_17_17_0_sva <= buf_acc_data_17_17_0_sva_mx0;
      buf_acc_data_17_17_45_1_sva <= buf_acc_data_17_17_45_1_sva_mx0;
      buf_acc_data_17_17_56_46_sva <= buf_acc_data_17_17_56_46_sva_mx0;
      buf_acc_data_0_0_0_sva <= buf_acc_data_0_0_0_sva_mx0;
      buf_acc_data_0_0_45_1_sva <= buf_acc_data_0_0_45_1_sva_mx0;
      buf_acc_data_0_0_56_46_sva <= buf_acc_data_0_0_56_46_sva_mx0;
      buf_acc_data_17_16_0_sva <= buf_acc_data_17_16_0_sva_mx0;
      buf_acc_data_17_16_45_1_sva <= buf_acc_data_17_16_45_1_sva_mx0;
      buf_acc_data_17_16_56_46_sva <= buf_acc_data_17_16_56_46_sva_mx0;
      buf_acc_data_0_1_0_sva <= buf_acc_data_0_1_0_sva_mx0;
      buf_acc_data_0_1_45_1_sva <= buf_acc_data_0_1_45_1_sva_mx0;
      buf_acc_data_0_1_56_46_sva <= buf_acc_data_0_1_56_46_sva_mx0;
      buf_acc_data_17_15_0_sva <= buf_acc_data_17_15_0_sva_mx0;
      buf_acc_data_17_15_45_1_sva <= buf_acc_data_17_15_45_1_sva_mx0;
      buf_acc_data_17_15_56_46_sva <= buf_acc_data_17_15_56_46_sva_mx0;
      buf_acc_data_0_2_0_sva <= buf_acc_data_0_2_0_sva_mx0;
      buf_acc_data_0_2_45_1_sva <= buf_acc_data_0_2_45_1_sva_mx0;
      buf_acc_data_0_2_56_46_sva <= buf_acc_data_0_2_56_46_sva_mx0;
      buf_acc_data_17_14_0_sva <= buf_acc_data_17_14_0_sva_mx0;
      buf_acc_data_17_14_45_1_sva <= buf_acc_data_17_14_45_1_sva_mx0;
      buf_acc_data_17_14_56_46_sva <= buf_acc_data_17_14_56_46_sva_mx0;
      buf_acc_data_0_3_0_sva <= buf_acc_data_0_3_0_sva_mx0;
      buf_acc_data_0_3_45_1_sva <= buf_acc_data_0_3_45_1_sva_mx0;
      buf_acc_data_0_3_56_46_sva <= buf_acc_data_0_3_56_46_sva_mx0;
      buf_acc_data_17_13_0_sva <= buf_acc_data_17_13_0_sva_mx0;
      buf_acc_data_17_13_45_1_sva <= buf_acc_data_17_13_45_1_sva_mx0;
      buf_acc_data_17_13_56_46_sva <= buf_acc_data_17_13_56_46_sva_mx0;
      buf_acc_data_0_4_0_sva <= buf_acc_data_0_4_0_sva_mx0;
      buf_acc_data_0_4_45_1_sva <= buf_acc_data_0_4_45_1_sva_mx0;
      buf_acc_data_0_4_56_46_sva <= buf_acc_data_0_4_56_46_sva_mx0;
      buf_acc_data_17_12_0_sva <= buf_acc_data_17_12_0_sva_mx0;
      buf_acc_data_17_12_45_1_sva <= buf_acc_data_17_12_45_1_sva_mx0;
      buf_acc_data_17_12_56_46_sva <= buf_acc_data_17_12_56_46_sva_mx0;
      buf_acc_data_0_5_0_sva <= buf_acc_data_0_5_0_sva_mx0;
      buf_acc_data_0_5_45_1_sva <= buf_acc_data_0_5_45_1_sva_mx0;
      buf_acc_data_0_5_56_46_sva <= buf_acc_data_0_5_56_46_sva_mx0;
      buf_acc_data_17_11_0_sva <= buf_acc_data_17_11_0_sva_mx0;
      buf_acc_data_17_11_45_1_sva <= buf_acc_data_17_11_45_1_sva_mx0;
      buf_acc_data_17_11_56_46_sva <= buf_acc_data_17_11_56_46_sva_mx0;
      buf_acc_data_0_6_0_sva <= buf_acc_data_0_6_0_sva_mx0;
      buf_acc_data_0_6_45_1_sva <= buf_acc_data_0_6_45_1_sva_mx0;
      buf_acc_data_0_6_56_46_sva <= buf_acc_data_0_6_56_46_sva_mx0;
      buf_acc_data_17_10_0_sva <= buf_acc_data_17_10_0_sva_mx0;
      buf_acc_data_17_10_45_1_sva <= buf_acc_data_17_10_45_1_sva_mx0;
      buf_acc_data_17_10_56_46_sva <= buf_acc_data_17_10_56_46_sva_mx0;
      buf_acc_data_0_7_0_sva <= buf_acc_data_0_7_0_sva_mx0;
      buf_acc_data_0_7_45_1_sva <= buf_acc_data_0_7_45_1_sva_mx0;
      buf_acc_data_0_7_56_46_sva <= buf_acc_data_0_7_56_46_sva_mx0;
      buf_acc_data_17_9_0_sva <= buf_acc_data_17_9_0_sva_mx0;
      buf_acc_data_17_9_45_1_sva <= buf_acc_data_17_9_45_1_sva_mx0;
      buf_acc_data_17_9_56_46_sva <= buf_acc_data_17_9_56_46_sva_mx0;
      buf_acc_data_0_8_0_sva <= buf_acc_data_0_8_0_sva_mx0;
      buf_acc_data_0_8_45_1_sva <= buf_acc_data_0_8_45_1_sva_mx0;
      buf_acc_data_0_8_56_46_sva <= buf_acc_data_0_8_56_46_sva_mx0;
      buf_acc_data_17_8_0_sva <= buf_acc_data_17_8_0_sva_mx0;
      buf_acc_data_17_8_45_1_sva <= buf_acc_data_17_8_45_1_sva_mx0;
      buf_acc_data_17_8_56_46_sva <= buf_acc_data_17_8_56_46_sva_mx0;
      buf_acc_data_0_9_0_sva <= buf_acc_data_0_9_0_sva_mx0;
      buf_acc_data_0_9_45_1_sva <= buf_acc_data_0_9_45_1_sva_mx0;
      buf_acc_data_0_9_56_46_sva <= buf_acc_data_0_9_56_46_sva_mx0;
      buf_acc_data_17_7_0_sva <= buf_acc_data_17_7_0_sva_mx0;
      buf_acc_data_17_7_45_1_sva <= buf_acc_data_17_7_45_1_sva_mx0;
      buf_acc_data_17_7_56_46_sva <= buf_acc_data_17_7_56_46_sva_mx0;
      buf_acc_data_0_10_0_sva <= buf_acc_data_0_10_0_sva_mx0;
      buf_acc_data_0_10_45_1_sva <= buf_acc_data_0_10_45_1_sva_mx0;
      buf_acc_data_0_10_56_46_sva <= buf_acc_data_0_10_56_46_sva_mx0;
      buf_acc_data_17_6_0_sva <= buf_acc_data_17_6_0_sva_mx0;
      buf_acc_data_17_6_45_1_sva <= buf_acc_data_17_6_45_1_sva_mx0;
      buf_acc_data_17_6_56_46_sva <= buf_acc_data_17_6_56_46_sva_mx0;
      buf_acc_data_0_11_0_sva <= buf_acc_data_0_11_0_sva_mx0;
      buf_acc_data_0_11_45_1_sva <= buf_acc_data_0_11_45_1_sva_mx0;
      buf_acc_data_0_11_56_46_sva <= buf_acc_data_0_11_56_46_sva_mx0;
      buf_acc_data_17_5_0_sva <= buf_acc_data_17_5_0_sva_mx0;
      buf_acc_data_17_5_45_1_sva <= buf_acc_data_17_5_45_1_sva_mx0;
      buf_acc_data_17_5_56_46_sva <= buf_acc_data_17_5_56_46_sva_mx0;
      buf_acc_data_0_12_0_sva <= buf_acc_data_0_12_0_sva_mx0;
      buf_acc_data_0_12_45_1_sva <= buf_acc_data_0_12_45_1_sva_mx0;
      buf_acc_data_0_12_56_46_sva <= buf_acc_data_0_12_56_46_sva_mx0;
      buf_acc_data_17_4_0_sva <= buf_acc_data_17_4_0_sva_mx0;
      buf_acc_data_17_4_45_1_sva <= buf_acc_data_17_4_45_1_sva_mx0;
      buf_acc_data_17_4_56_46_sva <= buf_acc_data_17_4_56_46_sva_mx0;
      buf_acc_data_0_13_0_sva <= buf_acc_data_0_13_0_sva_mx0;
      buf_acc_data_0_13_45_1_sva <= buf_acc_data_0_13_45_1_sva_mx0;
      buf_acc_data_0_13_56_46_sva <= buf_acc_data_0_13_56_46_sva_mx0;
      buf_acc_data_17_3_0_sva <= buf_acc_data_17_3_0_sva_mx0;
      buf_acc_data_17_3_45_1_sva <= buf_acc_data_17_3_45_1_sva_mx0;
      buf_acc_data_17_3_56_46_sva <= buf_acc_data_17_3_56_46_sva_mx0;
      buf_acc_data_0_14_0_sva <= buf_acc_data_0_14_0_sva_mx0;
      buf_acc_data_0_14_45_1_sva <= buf_acc_data_0_14_45_1_sva_mx0;
      buf_acc_data_0_14_56_46_sva <= buf_acc_data_0_14_56_46_sva_mx0;
      buf_acc_data_17_2_0_sva <= buf_acc_data_17_2_0_sva_mx0;
      buf_acc_data_17_2_45_1_sva <= buf_acc_data_17_2_45_1_sva_mx0;
      buf_acc_data_17_2_56_46_sva <= buf_acc_data_17_2_56_46_sva_mx0;
      buf_acc_data_0_15_0_sva <= buf_acc_data_0_15_0_sva_mx0;
      buf_acc_data_0_15_45_1_sva <= buf_acc_data_0_15_45_1_sva_mx0;
      buf_acc_data_0_15_56_46_sva <= buf_acc_data_0_15_56_46_sva_mx0;
      buf_acc_data_17_1_0_sva <= buf_acc_data_17_1_0_sva_mx0;
      buf_acc_data_17_1_45_1_sva <= buf_acc_data_17_1_45_1_sva_mx0;
      buf_acc_data_17_1_56_46_sva <= buf_acc_data_17_1_56_46_sva_mx0;
      buf_acc_data_0_16_0_sva <= buf_acc_data_0_16_0_sva_mx0;
      buf_acc_data_0_16_45_1_sva <= buf_acc_data_0_16_45_1_sva_mx0;
      buf_acc_data_0_16_56_46_sva <= buf_acc_data_0_16_56_46_sva_mx0;
      buf_acc_data_17_0_0_sva <= buf_acc_data_17_0_0_sva_mx0;
      buf_acc_data_17_0_45_1_sva <= buf_acc_data_17_0_45_1_sva_mx0;
      buf_acc_data_17_0_56_46_sva <= buf_acc_data_17_0_56_46_sva_mx0;
      buf_acc_data_0_17_0_sva <= buf_acc_data_0_17_0_sva_mx0;
      buf_acc_data_0_17_45_1_sva <= buf_acc_data_0_17_45_1_sva_mx0;
      buf_acc_data_0_17_56_46_sva <= buf_acc_data_0_17_56_46_sva_mx0;
      buf_acc_data_16_17_0_sva <= buf_acc_data_16_17_0_sva_mx0;
      buf_acc_data_16_17_45_1_sva <= buf_acc_data_16_17_45_1_sva_mx0;
      buf_acc_data_16_17_56_46_sva <= buf_acc_data_16_17_56_46_sva_mx0;
      buf_acc_data_1_0_0_sva <= buf_acc_data_1_0_0_sva_mx0;
      buf_acc_data_1_0_45_1_sva <= buf_acc_data_1_0_45_1_sva_mx0;
      buf_acc_data_1_0_56_46_sva <= buf_acc_data_1_0_56_46_sva_mx0;
      buf_acc_data_16_16_0_sva <= buf_acc_data_16_16_0_sva_mx0;
      buf_acc_data_16_16_45_1_sva <= buf_acc_data_16_16_45_1_sva_mx0;
      buf_acc_data_16_16_56_46_sva <= buf_acc_data_16_16_56_46_sva_mx0;
      buf_acc_data_1_1_0_sva <= buf_acc_data_1_1_0_sva_mx0;
      buf_acc_data_1_1_45_1_sva <= buf_acc_data_1_1_45_1_sva_mx0;
      buf_acc_data_1_1_56_46_sva <= buf_acc_data_1_1_56_46_sva_mx0;
      buf_acc_data_16_15_0_sva <= buf_acc_data_16_15_0_sva_mx0;
      buf_acc_data_16_15_45_1_sva <= buf_acc_data_16_15_45_1_sva_mx0;
      buf_acc_data_16_15_56_46_sva <= buf_acc_data_16_15_56_46_sva_mx0;
      buf_acc_data_1_2_0_sva <= buf_acc_data_1_2_0_sva_mx0;
      buf_acc_data_1_2_45_1_sva <= buf_acc_data_1_2_45_1_sva_mx0;
      buf_acc_data_1_2_56_46_sva <= buf_acc_data_1_2_56_46_sva_mx0;
      buf_acc_data_16_14_0_sva <= buf_acc_data_16_14_0_sva_mx0;
      buf_acc_data_16_14_45_1_sva <= buf_acc_data_16_14_45_1_sva_mx0;
      buf_acc_data_16_14_56_46_sva <= buf_acc_data_16_14_56_46_sva_mx0;
      buf_acc_data_1_3_0_sva <= buf_acc_data_1_3_0_sva_mx0;
      buf_acc_data_1_3_45_1_sva <= buf_acc_data_1_3_45_1_sva_mx0;
      buf_acc_data_1_3_56_46_sva <= buf_acc_data_1_3_56_46_sva_mx0;
      buf_acc_data_16_13_0_sva <= buf_acc_data_16_13_0_sva_mx0;
      buf_acc_data_16_13_45_1_sva <= buf_acc_data_16_13_45_1_sva_mx0;
      buf_acc_data_16_13_56_46_sva <= buf_acc_data_16_13_56_46_sva_mx0;
      buf_acc_data_1_4_0_sva <= buf_acc_data_1_4_0_sva_mx0;
      buf_acc_data_1_4_45_1_sva <= buf_acc_data_1_4_45_1_sva_mx0;
      buf_acc_data_1_4_56_46_sva <= buf_acc_data_1_4_56_46_sva_mx0;
      buf_acc_data_16_12_0_sva <= buf_acc_data_16_12_0_sva_mx0;
      buf_acc_data_16_12_45_1_sva <= buf_acc_data_16_12_45_1_sva_mx0;
      buf_acc_data_16_12_56_46_sva <= buf_acc_data_16_12_56_46_sva_mx0;
      buf_acc_data_1_5_0_sva <= buf_acc_data_1_5_0_sva_mx0;
      buf_acc_data_1_5_45_1_sva <= buf_acc_data_1_5_45_1_sva_mx0;
      buf_acc_data_1_5_56_46_sva <= buf_acc_data_1_5_56_46_sva_mx0;
      buf_acc_data_16_11_0_sva <= buf_acc_data_16_11_0_sva_mx0;
      buf_acc_data_16_11_45_1_sva <= buf_acc_data_16_11_45_1_sva_mx0;
      buf_acc_data_16_11_56_46_sva <= buf_acc_data_16_11_56_46_sva_mx0;
      buf_acc_data_1_6_0_sva <= buf_acc_data_1_6_0_sva_mx0;
      buf_acc_data_1_6_45_1_sva <= buf_acc_data_1_6_45_1_sva_mx0;
      buf_acc_data_1_6_56_46_sva <= buf_acc_data_1_6_56_46_sva_mx0;
      buf_acc_data_16_10_0_sva <= buf_acc_data_16_10_0_sva_mx0;
      buf_acc_data_16_10_45_1_sva <= buf_acc_data_16_10_45_1_sva_mx0;
      buf_acc_data_16_10_56_46_sva <= buf_acc_data_16_10_56_46_sva_mx0;
      buf_acc_data_1_7_0_sva <= buf_acc_data_1_7_0_sva_mx0;
      buf_acc_data_1_7_45_1_sva <= buf_acc_data_1_7_45_1_sva_mx0;
      buf_acc_data_1_7_56_46_sva <= buf_acc_data_1_7_56_46_sva_mx0;
      buf_acc_data_16_9_0_sva <= buf_acc_data_16_9_0_sva_mx0;
      buf_acc_data_16_9_45_1_sva <= buf_acc_data_16_9_45_1_sva_mx0;
      buf_acc_data_16_9_56_46_sva <= buf_acc_data_16_9_56_46_sva_mx0;
      buf_acc_data_1_8_0_sva <= buf_acc_data_1_8_0_sva_mx0;
      buf_acc_data_1_8_45_1_sva <= buf_acc_data_1_8_45_1_sva_mx0;
      buf_acc_data_1_8_56_46_sva <= buf_acc_data_1_8_56_46_sva_mx0;
      buf_acc_data_16_8_0_sva <= buf_acc_data_16_8_0_sva_mx0;
      buf_acc_data_16_8_45_1_sva <= buf_acc_data_16_8_45_1_sva_mx0;
      buf_acc_data_16_8_56_46_sva <= buf_acc_data_16_8_56_46_sva_mx0;
      buf_acc_data_1_9_0_sva <= buf_acc_data_1_9_0_sva_mx0;
      buf_acc_data_1_9_45_1_sva <= buf_acc_data_1_9_45_1_sva_mx0;
      buf_acc_data_1_9_56_46_sva <= buf_acc_data_1_9_56_46_sva_mx0;
      buf_acc_data_16_7_0_sva <= buf_acc_data_16_7_0_sva_mx0;
      buf_acc_data_16_7_45_1_sva <= buf_acc_data_16_7_45_1_sva_mx0;
      buf_acc_data_16_7_56_46_sva <= buf_acc_data_16_7_56_46_sva_mx0;
      buf_acc_data_1_10_0_sva <= buf_acc_data_1_10_0_sva_mx0;
      buf_acc_data_1_10_45_1_sva <= buf_acc_data_1_10_45_1_sva_mx0;
      buf_acc_data_1_10_56_46_sva <= buf_acc_data_1_10_56_46_sva_mx0;
      buf_acc_data_16_6_0_sva <= buf_acc_data_16_6_0_sva_mx0;
      buf_acc_data_16_6_45_1_sva <= buf_acc_data_16_6_45_1_sva_mx0;
      buf_acc_data_16_6_56_46_sva <= buf_acc_data_16_6_56_46_sva_mx0;
      buf_acc_data_1_11_0_sva <= buf_acc_data_1_11_0_sva_mx0;
      buf_acc_data_1_11_45_1_sva <= buf_acc_data_1_11_45_1_sva_mx0;
      buf_acc_data_1_11_56_46_sva <= buf_acc_data_1_11_56_46_sva_mx0;
      buf_acc_data_16_5_0_sva <= buf_acc_data_16_5_0_sva_mx0;
      buf_acc_data_16_5_45_1_sva <= buf_acc_data_16_5_45_1_sva_mx0;
      buf_acc_data_16_5_56_46_sva <= buf_acc_data_16_5_56_46_sva_mx0;
      buf_acc_data_1_12_0_sva <= buf_acc_data_1_12_0_sva_mx0;
      buf_acc_data_1_12_45_1_sva <= buf_acc_data_1_12_45_1_sva_mx0;
      buf_acc_data_1_12_56_46_sva <= buf_acc_data_1_12_56_46_sva_mx0;
      buf_acc_data_16_4_0_sva <= buf_acc_data_16_4_0_sva_mx0;
      buf_acc_data_16_4_45_1_sva <= buf_acc_data_16_4_45_1_sva_mx0;
      buf_acc_data_16_4_56_46_sva <= buf_acc_data_16_4_56_46_sva_mx0;
      buf_acc_data_1_13_0_sva <= buf_acc_data_1_13_0_sva_mx0;
      buf_acc_data_1_13_45_1_sva <= buf_acc_data_1_13_45_1_sva_mx0;
      buf_acc_data_1_13_56_46_sva <= buf_acc_data_1_13_56_46_sva_mx0;
      buf_acc_data_16_3_0_sva <= buf_acc_data_16_3_0_sva_mx0;
      buf_acc_data_16_3_45_1_sva <= buf_acc_data_16_3_45_1_sva_mx0;
      buf_acc_data_16_3_56_46_sva <= buf_acc_data_16_3_56_46_sva_mx0;
      buf_acc_data_1_14_0_sva <= buf_acc_data_1_14_0_sva_mx0;
      buf_acc_data_1_14_45_1_sva <= buf_acc_data_1_14_45_1_sva_mx0;
      buf_acc_data_1_14_56_46_sva <= buf_acc_data_1_14_56_46_sva_mx0;
      buf_acc_data_16_2_0_sva <= buf_acc_data_16_2_0_sva_mx0;
      buf_acc_data_16_2_45_1_sva <= buf_acc_data_16_2_45_1_sva_mx0;
      buf_acc_data_16_2_56_46_sva <= buf_acc_data_16_2_56_46_sva_mx0;
      buf_acc_data_1_15_0_sva <= buf_acc_data_1_15_0_sva_mx0;
      buf_acc_data_1_15_45_1_sva <= buf_acc_data_1_15_45_1_sva_mx0;
      buf_acc_data_1_15_56_46_sva <= buf_acc_data_1_15_56_46_sva_mx0;
      buf_acc_data_16_1_0_sva <= buf_acc_data_16_1_0_sva_mx0;
      buf_acc_data_16_1_45_1_sva <= buf_acc_data_16_1_45_1_sva_mx0;
      buf_acc_data_16_1_56_46_sva <= buf_acc_data_16_1_56_46_sva_mx0;
      buf_acc_data_1_16_0_sva <= buf_acc_data_1_16_0_sva_mx0;
      buf_acc_data_1_16_45_1_sva <= buf_acc_data_1_16_45_1_sva_mx0;
      buf_acc_data_1_16_56_46_sva <= buf_acc_data_1_16_56_46_sva_mx0;
      buf_acc_data_16_0_0_sva <= buf_acc_data_16_0_0_sva_mx0;
      buf_acc_data_16_0_45_1_sva <= buf_acc_data_16_0_45_1_sva_mx0;
      buf_acc_data_16_0_56_46_sva <= buf_acc_data_16_0_56_46_sva_mx0;
      buf_acc_data_1_17_0_sva <= buf_acc_data_1_17_0_sva_mx0;
      buf_acc_data_1_17_45_1_sva <= buf_acc_data_1_17_45_1_sva_mx0;
      buf_acc_data_1_17_56_46_sva <= buf_acc_data_1_17_56_46_sva_mx0;
      buf_acc_data_15_17_0_sva <= buf_acc_data_15_17_0_sva_mx0;
      buf_acc_data_15_17_45_1_sva <= buf_acc_data_15_17_45_1_sva_mx0;
      buf_acc_data_15_17_56_46_sva <= buf_acc_data_15_17_56_46_sva_mx0;
      buf_acc_data_2_0_0_sva <= buf_acc_data_2_0_0_sva_mx0;
      buf_acc_data_2_0_45_1_sva <= buf_acc_data_2_0_45_1_sva_mx0;
      buf_acc_data_2_0_56_46_sva <= buf_acc_data_2_0_56_46_sva_mx0;
      buf_acc_data_15_16_0_sva <= buf_acc_data_15_16_0_sva_mx0;
      buf_acc_data_15_16_45_1_sva <= buf_acc_data_15_16_45_1_sva_mx0;
      buf_acc_data_15_16_56_46_sva <= buf_acc_data_15_16_56_46_sva_mx0;
      buf_acc_data_2_1_0_sva <= buf_acc_data_2_1_0_sva_mx0;
      buf_acc_data_2_1_45_1_sva <= buf_acc_data_2_1_45_1_sva_mx0;
      buf_acc_data_2_1_56_46_sva <= buf_acc_data_2_1_56_46_sva_mx0;
      buf_acc_data_15_15_0_sva <= buf_acc_data_15_15_0_sva_mx0;
      buf_acc_data_15_15_45_1_sva <= buf_acc_data_15_15_45_1_sva_mx0;
      buf_acc_data_15_15_56_46_sva <= buf_acc_data_15_15_56_46_sva_mx0;
      buf_acc_data_2_2_0_sva <= buf_acc_data_2_2_0_sva_mx0;
      buf_acc_data_2_2_45_1_sva <= buf_acc_data_2_2_45_1_sva_mx0;
      buf_acc_data_2_2_56_46_sva <= buf_acc_data_2_2_56_46_sva_mx0;
      buf_acc_data_15_14_0_sva <= buf_acc_data_15_14_0_sva_mx0;
      buf_acc_data_15_14_45_1_sva <= buf_acc_data_15_14_45_1_sva_mx0;
      buf_acc_data_15_14_56_46_sva <= buf_acc_data_15_14_56_46_sva_mx0;
      buf_acc_data_2_3_0_sva <= buf_acc_data_2_3_0_sva_mx0;
      buf_acc_data_2_3_45_1_sva <= buf_acc_data_2_3_45_1_sva_mx0;
      buf_acc_data_2_3_56_46_sva <= buf_acc_data_2_3_56_46_sva_mx0;
      buf_acc_data_15_13_0_sva <= buf_acc_data_15_13_0_sva_mx0;
      buf_acc_data_15_13_45_1_sva <= buf_acc_data_15_13_45_1_sva_mx0;
      buf_acc_data_15_13_56_46_sva <= buf_acc_data_15_13_56_46_sva_mx0;
      buf_acc_data_2_4_0_sva <= buf_acc_data_2_4_0_sva_mx0;
      buf_acc_data_2_4_45_1_sva <= buf_acc_data_2_4_45_1_sva_mx0;
      buf_acc_data_2_4_56_46_sva <= buf_acc_data_2_4_56_46_sva_mx0;
      buf_acc_data_15_12_0_sva <= buf_acc_data_15_12_0_sva_mx0;
      buf_acc_data_15_12_45_1_sva <= buf_acc_data_15_12_45_1_sva_mx0;
      buf_acc_data_15_12_56_46_sva <= buf_acc_data_15_12_56_46_sva_mx0;
      buf_acc_data_2_5_0_sva <= buf_acc_data_2_5_0_sva_mx0;
      buf_acc_data_2_5_45_1_sva <= buf_acc_data_2_5_45_1_sva_mx0;
      buf_acc_data_2_5_56_46_sva <= buf_acc_data_2_5_56_46_sva_mx0;
      buf_acc_data_15_11_0_sva <= buf_acc_data_15_11_0_sva_mx0;
      buf_acc_data_15_11_45_1_sva <= buf_acc_data_15_11_45_1_sva_mx0;
      buf_acc_data_15_11_56_46_sva <= buf_acc_data_15_11_56_46_sva_mx0;
      buf_acc_data_2_6_0_sva <= buf_acc_data_2_6_0_sva_mx0;
      buf_acc_data_2_6_45_1_sva <= buf_acc_data_2_6_45_1_sva_mx0;
      buf_acc_data_2_6_56_46_sva <= buf_acc_data_2_6_56_46_sva_mx0;
      buf_acc_data_15_10_0_sva <= buf_acc_data_15_10_0_sva_mx0;
      buf_acc_data_15_10_45_1_sva <= buf_acc_data_15_10_45_1_sva_mx0;
      buf_acc_data_15_10_56_46_sva <= buf_acc_data_15_10_56_46_sva_mx0;
      buf_acc_data_2_7_0_sva <= buf_acc_data_2_7_0_sva_mx0;
      buf_acc_data_2_7_45_1_sva <= buf_acc_data_2_7_45_1_sva_mx0;
      buf_acc_data_2_7_56_46_sva <= buf_acc_data_2_7_56_46_sva_mx0;
      buf_acc_data_15_9_0_sva <= buf_acc_data_15_9_0_sva_mx0;
      buf_acc_data_15_9_45_1_sva <= buf_acc_data_15_9_45_1_sva_mx0;
      buf_acc_data_15_9_56_46_sva <= buf_acc_data_15_9_56_46_sva_mx0;
      buf_acc_data_2_8_0_sva <= buf_acc_data_2_8_0_sva_mx0;
      buf_acc_data_2_8_45_1_sva <= buf_acc_data_2_8_45_1_sva_mx0;
      buf_acc_data_2_8_56_46_sva <= buf_acc_data_2_8_56_46_sva_mx0;
      buf_acc_data_15_8_0_sva <= buf_acc_data_15_8_0_sva_mx0;
      buf_acc_data_15_8_45_1_sva <= buf_acc_data_15_8_45_1_sva_mx0;
      buf_acc_data_15_8_56_46_sva <= buf_acc_data_15_8_56_46_sva_mx0;
      buf_acc_data_2_9_0_sva <= buf_acc_data_2_9_0_sva_mx0;
      buf_acc_data_2_9_45_1_sva <= buf_acc_data_2_9_45_1_sva_mx0;
      buf_acc_data_2_9_56_46_sva <= buf_acc_data_2_9_56_46_sva_mx0;
      buf_acc_data_15_7_0_sva <= buf_acc_data_15_7_0_sva_mx0;
      buf_acc_data_15_7_45_1_sva <= buf_acc_data_15_7_45_1_sva_mx0;
      buf_acc_data_15_7_56_46_sva <= buf_acc_data_15_7_56_46_sva_mx0;
      buf_acc_data_2_10_0_sva <= buf_acc_data_2_10_0_sva_mx0;
      buf_acc_data_2_10_45_1_sva <= buf_acc_data_2_10_45_1_sva_mx0;
      buf_acc_data_2_10_56_46_sva <= buf_acc_data_2_10_56_46_sva_mx0;
      buf_acc_data_15_6_0_sva <= buf_acc_data_15_6_0_sva_mx0;
      buf_acc_data_15_6_45_1_sva <= buf_acc_data_15_6_45_1_sva_mx0;
      buf_acc_data_15_6_56_46_sva <= buf_acc_data_15_6_56_46_sva_mx0;
      buf_acc_data_2_11_0_sva <= buf_acc_data_2_11_0_sva_mx0;
      buf_acc_data_2_11_45_1_sva <= buf_acc_data_2_11_45_1_sva_mx0;
      buf_acc_data_2_11_56_46_sva <= buf_acc_data_2_11_56_46_sva_mx0;
      buf_acc_data_15_5_0_sva <= buf_acc_data_15_5_0_sva_mx0;
      buf_acc_data_15_5_45_1_sva <= buf_acc_data_15_5_45_1_sva_mx0;
      buf_acc_data_15_5_56_46_sva <= buf_acc_data_15_5_56_46_sva_mx0;
      buf_acc_data_2_12_0_sva <= buf_acc_data_2_12_0_sva_mx0;
      buf_acc_data_2_12_45_1_sva <= buf_acc_data_2_12_45_1_sva_mx0;
      buf_acc_data_2_12_56_46_sva <= buf_acc_data_2_12_56_46_sva_mx0;
      buf_acc_data_15_4_0_sva <= buf_acc_data_15_4_0_sva_mx0;
      buf_acc_data_15_4_45_1_sva <= buf_acc_data_15_4_45_1_sva_mx0;
      buf_acc_data_15_4_56_46_sva <= buf_acc_data_15_4_56_46_sva_mx0;
      buf_acc_data_2_13_0_sva <= buf_acc_data_2_13_0_sva_mx0;
      buf_acc_data_2_13_45_1_sva <= buf_acc_data_2_13_45_1_sva_mx0;
      buf_acc_data_2_13_56_46_sva <= buf_acc_data_2_13_56_46_sva_mx0;
      buf_acc_data_15_3_0_sva <= buf_acc_data_15_3_0_sva_mx0;
      buf_acc_data_15_3_45_1_sva <= buf_acc_data_15_3_45_1_sva_mx0;
      buf_acc_data_15_3_56_46_sva <= buf_acc_data_15_3_56_46_sva_mx0;
      buf_acc_data_2_14_0_sva <= buf_acc_data_2_14_0_sva_mx0;
      buf_acc_data_2_14_45_1_sva <= buf_acc_data_2_14_45_1_sva_mx0;
      buf_acc_data_2_14_56_46_sva <= buf_acc_data_2_14_56_46_sva_mx0;
      buf_acc_data_15_2_0_sva <= buf_acc_data_15_2_0_sva_mx0;
      buf_acc_data_15_2_45_1_sva <= buf_acc_data_15_2_45_1_sva_mx0;
      buf_acc_data_15_2_56_46_sva <= buf_acc_data_15_2_56_46_sva_mx0;
      buf_acc_data_2_15_0_sva <= buf_acc_data_2_15_0_sva_mx0;
      buf_acc_data_2_15_45_1_sva <= buf_acc_data_2_15_45_1_sva_mx0;
      buf_acc_data_2_15_56_46_sva <= buf_acc_data_2_15_56_46_sva_mx0;
      buf_acc_data_15_1_0_sva <= buf_acc_data_15_1_0_sva_mx0;
      buf_acc_data_15_1_45_1_sva <= buf_acc_data_15_1_45_1_sva_mx0;
      buf_acc_data_15_1_56_46_sva <= buf_acc_data_15_1_56_46_sva_mx0;
      buf_acc_data_2_16_0_sva <= buf_acc_data_2_16_0_sva_mx0;
      buf_acc_data_2_16_45_1_sva <= buf_acc_data_2_16_45_1_sva_mx0;
      buf_acc_data_2_16_56_46_sva <= buf_acc_data_2_16_56_46_sva_mx0;
      buf_acc_data_15_0_0_sva <= buf_acc_data_15_0_0_sva_mx0;
      buf_acc_data_15_0_45_1_sva <= buf_acc_data_15_0_45_1_sva_mx0;
      buf_acc_data_15_0_56_46_sva <= buf_acc_data_15_0_56_46_sva_mx0;
      buf_acc_data_2_17_0_sva <= buf_acc_data_2_17_0_sva_mx0;
      buf_acc_data_2_17_45_1_sva <= buf_acc_data_2_17_45_1_sva_mx0;
      buf_acc_data_2_17_56_46_sva <= buf_acc_data_2_17_56_46_sva_mx0;
      buf_acc_data_14_17_0_sva <= buf_acc_data_14_17_0_sva_mx0;
      buf_acc_data_14_17_45_1_sva <= buf_acc_data_14_17_45_1_sva_mx0;
      buf_acc_data_14_17_56_46_sva <= buf_acc_data_14_17_56_46_sva_mx0;
      buf_acc_data_3_0_0_sva <= buf_acc_data_3_0_0_sva_mx0;
      buf_acc_data_3_0_45_1_sva <= buf_acc_data_3_0_45_1_sva_mx0;
      buf_acc_data_3_0_56_46_sva <= buf_acc_data_3_0_56_46_sva_mx0;
      buf_acc_data_14_16_0_sva <= buf_acc_data_14_16_0_sva_mx0;
      buf_acc_data_14_16_45_1_sva <= buf_acc_data_14_16_45_1_sva_mx0;
      buf_acc_data_14_16_56_46_sva <= buf_acc_data_14_16_56_46_sva_mx0;
      buf_acc_data_3_1_0_sva <= buf_acc_data_3_1_0_sva_mx0;
      buf_acc_data_3_1_45_1_sva <= buf_acc_data_3_1_45_1_sva_mx0;
      buf_acc_data_3_1_56_46_sva <= buf_acc_data_3_1_56_46_sva_mx0;
      buf_acc_data_14_15_0_sva <= buf_acc_data_14_15_0_sva_mx0;
      buf_acc_data_14_15_45_1_sva <= buf_acc_data_14_15_45_1_sva_mx0;
      buf_acc_data_14_15_56_46_sva <= buf_acc_data_14_15_56_46_sva_mx0;
      buf_acc_data_3_2_0_sva <= buf_acc_data_3_2_0_sva_mx0;
      buf_acc_data_3_2_45_1_sva <= buf_acc_data_3_2_45_1_sva_mx0;
      buf_acc_data_3_2_56_46_sva <= buf_acc_data_3_2_56_46_sva_mx0;
      buf_acc_data_14_14_0_sva <= buf_acc_data_14_14_0_sva_mx0;
      buf_acc_data_14_14_45_1_sva <= buf_acc_data_14_14_45_1_sva_mx0;
      buf_acc_data_14_14_56_46_sva <= buf_acc_data_14_14_56_46_sva_mx0;
      buf_acc_data_3_3_0_sva <= buf_acc_data_3_3_0_sva_mx0;
      buf_acc_data_3_3_45_1_sva <= buf_acc_data_3_3_45_1_sva_mx0;
      buf_acc_data_3_3_56_46_sva <= buf_acc_data_3_3_56_46_sva_mx0;
      buf_acc_data_14_13_0_sva <= buf_acc_data_14_13_0_sva_mx0;
      buf_acc_data_14_13_45_1_sva <= buf_acc_data_14_13_45_1_sva_mx0;
      buf_acc_data_14_13_56_46_sva <= buf_acc_data_14_13_56_46_sva_mx0;
      buf_acc_data_3_4_0_sva <= buf_acc_data_3_4_0_sva_mx0;
      buf_acc_data_3_4_45_1_sva <= buf_acc_data_3_4_45_1_sva_mx0;
      buf_acc_data_3_4_56_46_sva <= buf_acc_data_3_4_56_46_sva_mx0;
      buf_acc_data_14_12_0_sva <= buf_acc_data_14_12_0_sva_mx0;
      buf_acc_data_14_12_45_1_sva <= buf_acc_data_14_12_45_1_sva_mx0;
      buf_acc_data_14_12_56_46_sva <= buf_acc_data_14_12_56_46_sva_mx0;
      buf_acc_data_3_5_0_sva <= buf_acc_data_3_5_0_sva_mx0;
      buf_acc_data_3_5_45_1_sva <= buf_acc_data_3_5_45_1_sva_mx0;
      buf_acc_data_3_5_56_46_sva <= buf_acc_data_3_5_56_46_sva_mx0;
      buf_acc_data_14_11_0_sva <= buf_acc_data_14_11_0_sva_mx0;
      buf_acc_data_14_11_45_1_sva <= buf_acc_data_14_11_45_1_sva_mx0;
      buf_acc_data_14_11_56_46_sva <= buf_acc_data_14_11_56_46_sva_mx0;
      buf_acc_data_3_6_0_sva <= buf_acc_data_3_6_0_sva_mx0;
      buf_acc_data_3_6_45_1_sva <= buf_acc_data_3_6_45_1_sva_mx0;
      buf_acc_data_3_6_56_46_sva <= buf_acc_data_3_6_56_46_sva_mx0;
      buf_acc_data_14_10_0_sva <= buf_acc_data_14_10_0_sva_mx0;
      buf_acc_data_14_10_45_1_sva <= buf_acc_data_14_10_45_1_sva_mx0;
      buf_acc_data_14_10_56_46_sva <= buf_acc_data_14_10_56_46_sva_mx0;
      buf_acc_data_3_7_0_sva <= buf_acc_data_3_7_0_sva_mx0;
      buf_acc_data_3_7_45_1_sva <= buf_acc_data_3_7_45_1_sva_mx0;
      buf_acc_data_3_7_56_46_sva <= buf_acc_data_3_7_56_46_sva_mx0;
      buf_acc_data_14_9_0_sva <= buf_acc_data_14_9_0_sva_mx0;
      buf_acc_data_14_9_45_1_sva <= buf_acc_data_14_9_45_1_sva_mx0;
      buf_acc_data_14_9_56_46_sva <= buf_acc_data_14_9_56_46_sva_mx0;
      buf_acc_data_3_8_0_sva <= buf_acc_data_3_8_0_sva_mx0;
      buf_acc_data_3_8_45_1_sva <= buf_acc_data_3_8_45_1_sva_mx0;
      buf_acc_data_3_8_56_46_sva <= buf_acc_data_3_8_56_46_sva_mx0;
      buf_acc_data_14_8_0_sva <= buf_acc_data_14_8_0_sva_mx0;
      buf_acc_data_14_8_45_1_sva <= buf_acc_data_14_8_45_1_sva_mx0;
      buf_acc_data_14_8_56_46_sva <= buf_acc_data_14_8_56_46_sva_mx0;
      buf_acc_data_3_9_0_sva <= buf_acc_data_3_9_0_sva_mx0;
      buf_acc_data_3_9_45_1_sva <= buf_acc_data_3_9_45_1_sva_mx0;
      buf_acc_data_3_9_56_46_sva <= buf_acc_data_3_9_56_46_sva_mx0;
      buf_acc_data_14_7_0_sva <= buf_acc_data_14_7_0_sva_mx0;
      buf_acc_data_14_7_45_1_sva <= buf_acc_data_14_7_45_1_sva_mx0;
      buf_acc_data_14_7_56_46_sva <= buf_acc_data_14_7_56_46_sva_mx0;
      buf_acc_data_3_10_0_sva <= buf_acc_data_3_10_0_sva_mx0;
      buf_acc_data_3_10_45_1_sva <= buf_acc_data_3_10_45_1_sva_mx0;
      buf_acc_data_3_10_56_46_sva <= buf_acc_data_3_10_56_46_sva_mx0;
      buf_acc_data_14_6_0_sva <= buf_acc_data_14_6_0_sva_mx0;
      buf_acc_data_14_6_45_1_sva <= buf_acc_data_14_6_45_1_sva_mx0;
      buf_acc_data_14_6_56_46_sva <= buf_acc_data_14_6_56_46_sva_mx0;
      buf_acc_data_3_11_0_sva <= buf_acc_data_3_11_0_sva_mx0;
      buf_acc_data_3_11_45_1_sva <= buf_acc_data_3_11_45_1_sva_mx0;
      buf_acc_data_3_11_56_46_sva <= buf_acc_data_3_11_56_46_sva_mx0;
      buf_acc_data_14_5_0_sva <= buf_acc_data_14_5_0_sva_mx0;
      buf_acc_data_14_5_45_1_sva <= buf_acc_data_14_5_45_1_sva_mx0;
      buf_acc_data_14_5_56_46_sva <= buf_acc_data_14_5_56_46_sva_mx0;
      buf_acc_data_3_12_0_sva <= buf_acc_data_3_12_0_sva_mx0;
      buf_acc_data_3_12_45_1_sva <= buf_acc_data_3_12_45_1_sva_mx0;
      buf_acc_data_3_12_56_46_sva <= buf_acc_data_3_12_56_46_sva_mx0;
      buf_acc_data_14_4_0_sva <= buf_acc_data_14_4_0_sva_mx0;
      buf_acc_data_14_4_45_1_sva <= buf_acc_data_14_4_45_1_sva_mx0;
      buf_acc_data_14_4_56_46_sva <= buf_acc_data_14_4_56_46_sva_mx0;
      buf_acc_data_3_13_0_sva <= buf_acc_data_3_13_0_sva_mx0;
      buf_acc_data_3_13_45_1_sva <= buf_acc_data_3_13_45_1_sva_mx0;
      buf_acc_data_3_13_56_46_sva <= buf_acc_data_3_13_56_46_sva_mx0;
      buf_acc_data_14_3_0_sva <= buf_acc_data_14_3_0_sva_mx0;
      buf_acc_data_14_3_45_1_sva <= buf_acc_data_14_3_45_1_sva_mx0;
      buf_acc_data_14_3_56_46_sva <= buf_acc_data_14_3_56_46_sva_mx0;
      buf_acc_data_3_14_0_sva <= buf_acc_data_3_14_0_sva_mx0;
      buf_acc_data_3_14_45_1_sva <= buf_acc_data_3_14_45_1_sva_mx0;
      buf_acc_data_3_14_56_46_sva <= buf_acc_data_3_14_56_46_sva_mx0;
      buf_acc_data_14_2_0_sva <= buf_acc_data_14_2_0_sva_mx0;
      buf_acc_data_14_2_45_1_sva <= buf_acc_data_14_2_45_1_sva_mx0;
      buf_acc_data_14_2_56_46_sva <= buf_acc_data_14_2_56_46_sva_mx0;
      buf_acc_data_3_15_0_sva <= buf_acc_data_3_15_0_sva_mx0;
      buf_acc_data_3_15_45_1_sva <= buf_acc_data_3_15_45_1_sva_mx0;
      buf_acc_data_3_15_56_46_sva <= buf_acc_data_3_15_56_46_sva_mx0;
      buf_acc_data_14_1_0_sva <= buf_acc_data_14_1_0_sva_mx0;
      buf_acc_data_14_1_45_1_sva <= buf_acc_data_14_1_45_1_sva_mx0;
      buf_acc_data_14_1_56_46_sva <= buf_acc_data_14_1_56_46_sva_mx0;
      buf_acc_data_3_16_0_sva <= buf_acc_data_3_16_0_sva_mx0;
      buf_acc_data_3_16_45_1_sva <= buf_acc_data_3_16_45_1_sva_mx0;
      buf_acc_data_3_16_56_46_sva <= buf_acc_data_3_16_56_46_sva_mx0;
      buf_acc_data_14_0_0_sva <= buf_acc_data_14_0_0_sva_mx0;
      buf_acc_data_14_0_45_1_sva <= buf_acc_data_14_0_45_1_sva_mx0;
      buf_acc_data_14_0_56_46_sva <= buf_acc_data_14_0_56_46_sva_mx0;
      buf_acc_data_3_17_0_sva <= buf_acc_data_3_17_0_sva_mx0;
      buf_acc_data_3_17_45_1_sva <= buf_acc_data_3_17_45_1_sva_mx0;
      buf_acc_data_3_17_56_46_sva <= buf_acc_data_3_17_56_46_sva_mx0;
      buf_acc_data_13_17_0_sva <= buf_acc_data_13_17_0_sva_mx0;
      buf_acc_data_13_17_45_1_sva <= buf_acc_data_13_17_45_1_sva_mx0;
      buf_acc_data_13_17_56_46_sva <= buf_acc_data_13_17_56_46_sva_mx0;
      buf_acc_data_4_0_0_sva <= buf_acc_data_4_0_0_sva_mx0;
      buf_acc_data_4_0_45_1_sva <= buf_acc_data_4_0_45_1_sva_mx0;
      buf_acc_data_4_0_56_46_sva <= buf_acc_data_4_0_56_46_sva_mx0;
      buf_acc_data_13_16_0_sva <= buf_acc_data_13_16_0_sva_mx0;
      buf_acc_data_13_16_45_1_sva <= buf_acc_data_13_16_45_1_sva_mx0;
      buf_acc_data_13_16_56_46_sva <= buf_acc_data_13_16_56_46_sva_mx0;
      buf_acc_data_4_1_0_sva <= buf_acc_data_4_1_0_sva_mx0;
      buf_acc_data_4_1_45_1_sva <= buf_acc_data_4_1_45_1_sva_mx0;
      buf_acc_data_4_1_56_46_sva <= buf_acc_data_4_1_56_46_sva_mx0;
      buf_acc_data_13_15_0_sva <= buf_acc_data_13_15_0_sva_mx0;
      buf_acc_data_13_15_45_1_sva <= buf_acc_data_13_15_45_1_sva_mx0;
      buf_acc_data_13_15_56_46_sva <= buf_acc_data_13_15_56_46_sva_mx0;
      buf_acc_data_4_2_0_sva <= buf_acc_data_4_2_0_sva_mx0;
      buf_acc_data_4_2_45_1_sva <= buf_acc_data_4_2_45_1_sva_mx0;
      buf_acc_data_4_2_56_46_sva <= buf_acc_data_4_2_56_46_sva_mx0;
      buf_acc_data_13_14_0_sva <= buf_acc_data_13_14_0_sva_mx0;
      buf_acc_data_13_14_45_1_sva <= buf_acc_data_13_14_45_1_sva_mx0;
      buf_acc_data_13_14_56_46_sva <= buf_acc_data_13_14_56_46_sva_mx0;
      buf_acc_data_4_3_0_sva <= buf_acc_data_4_3_0_sva_mx0;
      buf_acc_data_4_3_45_1_sva <= buf_acc_data_4_3_45_1_sva_mx0;
      buf_acc_data_4_3_56_46_sva <= buf_acc_data_4_3_56_46_sva_mx0;
      buf_acc_data_13_13_0_sva <= buf_acc_data_13_13_0_sva_mx0;
      buf_acc_data_13_13_45_1_sva <= buf_acc_data_13_13_45_1_sva_mx0;
      buf_acc_data_13_13_56_46_sva <= buf_acc_data_13_13_56_46_sva_mx0;
      buf_acc_data_4_4_0_sva <= buf_acc_data_4_4_0_sva_mx0;
      buf_acc_data_4_4_45_1_sva <= buf_acc_data_4_4_45_1_sva_mx0;
      buf_acc_data_4_4_56_46_sva <= buf_acc_data_4_4_56_46_sva_mx0;
      buf_acc_data_13_12_0_sva <= buf_acc_data_13_12_0_sva_mx0;
      buf_acc_data_13_12_45_1_sva <= buf_acc_data_13_12_45_1_sva_mx0;
      buf_acc_data_13_12_56_46_sva <= buf_acc_data_13_12_56_46_sva_mx0;
      buf_acc_data_4_5_0_sva <= buf_acc_data_4_5_0_sva_mx0;
      buf_acc_data_4_5_45_1_sva <= buf_acc_data_4_5_45_1_sva_mx0;
      buf_acc_data_4_5_56_46_sva <= buf_acc_data_4_5_56_46_sva_mx0;
      buf_acc_data_13_11_0_sva <= buf_acc_data_13_11_0_sva_mx0;
      buf_acc_data_13_11_45_1_sva <= buf_acc_data_13_11_45_1_sva_mx0;
      buf_acc_data_13_11_56_46_sva <= buf_acc_data_13_11_56_46_sva_mx0;
      buf_acc_data_4_6_0_sva <= buf_acc_data_4_6_0_sva_mx0;
      buf_acc_data_4_6_45_1_sva <= buf_acc_data_4_6_45_1_sva_mx0;
      buf_acc_data_4_6_56_46_sva <= buf_acc_data_4_6_56_46_sva_mx0;
      buf_acc_data_13_10_0_sva <= buf_acc_data_13_10_0_sva_mx0;
      buf_acc_data_13_10_45_1_sva <= buf_acc_data_13_10_45_1_sva_mx0;
      buf_acc_data_13_10_56_46_sva <= buf_acc_data_13_10_56_46_sva_mx0;
      buf_acc_data_4_7_0_sva <= buf_acc_data_4_7_0_sva_mx0;
      buf_acc_data_4_7_45_1_sva <= buf_acc_data_4_7_45_1_sva_mx0;
      buf_acc_data_4_7_56_46_sva <= buf_acc_data_4_7_56_46_sva_mx0;
      buf_acc_data_13_9_0_sva <= buf_acc_data_13_9_0_sva_mx0;
      buf_acc_data_13_9_45_1_sva <= buf_acc_data_13_9_45_1_sva_mx0;
      buf_acc_data_13_9_56_46_sva <= buf_acc_data_13_9_56_46_sva_mx0;
      buf_acc_data_4_8_0_sva <= buf_acc_data_4_8_0_sva_mx0;
      buf_acc_data_4_8_45_1_sva <= buf_acc_data_4_8_45_1_sva_mx0;
      buf_acc_data_4_8_56_46_sva <= buf_acc_data_4_8_56_46_sva_mx0;
      buf_acc_data_13_8_0_sva <= buf_acc_data_13_8_0_sva_mx0;
      buf_acc_data_13_8_45_1_sva <= buf_acc_data_13_8_45_1_sva_mx0;
      buf_acc_data_13_8_56_46_sva <= buf_acc_data_13_8_56_46_sva_mx0;
      buf_acc_data_4_9_0_sva <= buf_acc_data_4_9_0_sva_mx0;
      buf_acc_data_4_9_45_1_sva <= buf_acc_data_4_9_45_1_sva_mx0;
      buf_acc_data_4_9_56_46_sva <= buf_acc_data_4_9_56_46_sva_mx0;
      buf_acc_data_13_7_0_sva <= buf_acc_data_13_7_0_sva_mx0;
      buf_acc_data_13_7_45_1_sva <= buf_acc_data_13_7_45_1_sva_mx0;
      buf_acc_data_13_7_56_46_sva <= buf_acc_data_13_7_56_46_sva_mx0;
      buf_acc_data_4_10_0_sva <= buf_acc_data_4_10_0_sva_mx0;
      buf_acc_data_4_10_45_1_sva <= buf_acc_data_4_10_45_1_sva_mx0;
      buf_acc_data_4_10_56_46_sva <= buf_acc_data_4_10_56_46_sva_mx0;
      buf_acc_data_13_6_0_sva <= buf_acc_data_13_6_0_sva_mx0;
      buf_acc_data_13_6_45_1_sva <= buf_acc_data_13_6_45_1_sva_mx0;
      buf_acc_data_13_6_56_46_sva <= buf_acc_data_13_6_56_46_sva_mx0;
      buf_acc_data_4_11_0_sva <= buf_acc_data_4_11_0_sva_mx0;
      buf_acc_data_4_11_45_1_sva <= buf_acc_data_4_11_45_1_sva_mx0;
      buf_acc_data_4_11_56_46_sva <= buf_acc_data_4_11_56_46_sva_mx0;
      buf_acc_data_13_5_0_sva <= buf_acc_data_13_5_0_sva_mx0;
      buf_acc_data_13_5_45_1_sva <= buf_acc_data_13_5_45_1_sva_mx0;
      buf_acc_data_13_5_56_46_sva <= buf_acc_data_13_5_56_46_sva_mx0;
      buf_acc_data_4_12_0_sva <= buf_acc_data_4_12_0_sva_mx0;
      buf_acc_data_4_12_45_1_sva <= buf_acc_data_4_12_45_1_sva_mx0;
      buf_acc_data_4_12_56_46_sva <= buf_acc_data_4_12_56_46_sva_mx0;
      buf_acc_data_13_4_0_sva <= buf_acc_data_13_4_0_sva_mx0;
      buf_acc_data_13_4_45_1_sva <= buf_acc_data_13_4_45_1_sva_mx0;
      buf_acc_data_13_4_56_46_sva <= buf_acc_data_13_4_56_46_sva_mx0;
      buf_acc_data_4_13_0_sva <= buf_acc_data_4_13_0_sva_mx0;
      buf_acc_data_4_13_45_1_sva <= buf_acc_data_4_13_45_1_sva_mx0;
      buf_acc_data_4_13_56_46_sva <= buf_acc_data_4_13_56_46_sva_mx0;
      buf_acc_data_13_3_0_sva <= buf_acc_data_13_3_0_sva_mx0;
      buf_acc_data_13_3_45_1_sva <= buf_acc_data_13_3_45_1_sva_mx0;
      buf_acc_data_13_3_56_46_sva <= buf_acc_data_13_3_56_46_sva_mx0;
      buf_acc_data_4_14_0_sva <= buf_acc_data_4_14_0_sva_mx0;
      buf_acc_data_4_14_45_1_sva <= buf_acc_data_4_14_45_1_sva_mx0;
      buf_acc_data_4_14_56_46_sva <= buf_acc_data_4_14_56_46_sva_mx0;
      buf_acc_data_13_2_0_sva <= buf_acc_data_13_2_0_sva_mx0;
      buf_acc_data_13_2_45_1_sva <= buf_acc_data_13_2_45_1_sva_mx0;
      buf_acc_data_13_2_56_46_sva <= buf_acc_data_13_2_56_46_sva_mx0;
      buf_acc_data_4_15_0_sva <= buf_acc_data_4_15_0_sva_mx0;
      buf_acc_data_4_15_45_1_sva <= buf_acc_data_4_15_45_1_sva_mx0;
      buf_acc_data_4_15_56_46_sva <= buf_acc_data_4_15_56_46_sva_mx0;
      buf_acc_data_13_1_0_sva <= buf_acc_data_13_1_0_sva_mx0;
      buf_acc_data_13_1_45_1_sva <= buf_acc_data_13_1_45_1_sva_mx0;
      buf_acc_data_13_1_56_46_sva <= buf_acc_data_13_1_56_46_sva_mx0;
      buf_acc_data_4_16_0_sva <= buf_acc_data_4_16_0_sva_mx0;
      buf_acc_data_4_16_45_1_sva <= buf_acc_data_4_16_45_1_sva_mx0;
      buf_acc_data_4_16_56_46_sva <= buf_acc_data_4_16_56_46_sva_mx0;
      buf_acc_data_13_0_0_sva <= buf_acc_data_13_0_0_sva_mx0;
      buf_acc_data_13_0_45_1_sva <= buf_acc_data_13_0_45_1_sva_mx0;
      buf_acc_data_13_0_56_46_sva <= buf_acc_data_13_0_56_46_sva_mx0;
      buf_acc_data_4_17_0_sva <= buf_acc_data_4_17_0_sva_mx0;
      buf_acc_data_4_17_45_1_sva <= buf_acc_data_4_17_45_1_sva_mx0;
      buf_acc_data_4_17_56_46_sva <= buf_acc_data_4_17_56_46_sva_mx0;
      buf_acc_data_12_17_0_sva <= buf_acc_data_12_17_0_sva_mx0;
      buf_acc_data_12_17_45_1_sva <= buf_acc_data_12_17_45_1_sva_mx0;
      buf_acc_data_12_17_56_46_sva <= buf_acc_data_12_17_56_46_sva_mx0;
      buf_acc_data_5_0_0_sva <= buf_acc_data_5_0_0_sva_mx0;
      buf_acc_data_5_0_45_1_sva <= buf_acc_data_5_0_45_1_sva_mx0;
      buf_acc_data_5_0_56_46_sva <= buf_acc_data_5_0_56_46_sva_mx0;
      buf_acc_data_12_16_0_sva <= buf_acc_data_12_16_0_sva_mx0;
      buf_acc_data_12_16_45_1_sva <= buf_acc_data_12_16_45_1_sva_mx0;
      buf_acc_data_12_16_56_46_sva <= buf_acc_data_12_16_56_46_sva_mx0;
      buf_acc_data_5_1_0_sva <= buf_acc_data_5_1_0_sva_mx0;
      buf_acc_data_5_1_45_1_sva <= buf_acc_data_5_1_45_1_sva_mx0;
      buf_acc_data_5_1_56_46_sva <= buf_acc_data_5_1_56_46_sva_mx0;
      buf_acc_data_12_15_0_sva <= buf_acc_data_12_15_0_sva_mx0;
      buf_acc_data_12_15_45_1_sva <= buf_acc_data_12_15_45_1_sva_mx0;
      buf_acc_data_12_15_56_46_sva <= buf_acc_data_12_15_56_46_sva_mx0;
      buf_acc_data_5_2_0_sva <= buf_acc_data_5_2_0_sva_mx0;
      buf_acc_data_5_2_45_1_sva <= buf_acc_data_5_2_45_1_sva_mx0;
      buf_acc_data_5_2_56_46_sva <= buf_acc_data_5_2_56_46_sva_mx0;
      buf_acc_data_12_14_0_sva <= buf_acc_data_12_14_0_sva_mx0;
      buf_acc_data_12_14_45_1_sva <= buf_acc_data_12_14_45_1_sva_mx0;
      buf_acc_data_12_14_56_46_sva <= buf_acc_data_12_14_56_46_sva_mx0;
      buf_acc_data_5_3_0_sva <= buf_acc_data_5_3_0_sva_mx0;
      buf_acc_data_5_3_45_1_sva <= buf_acc_data_5_3_45_1_sva_mx0;
      buf_acc_data_5_3_56_46_sva <= buf_acc_data_5_3_56_46_sva_mx0;
      buf_acc_data_12_13_0_sva <= buf_acc_data_12_13_0_sva_mx0;
      buf_acc_data_12_13_45_1_sva <= buf_acc_data_12_13_45_1_sva_mx0;
      buf_acc_data_12_13_56_46_sva <= buf_acc_data_12_13_56_46_sva_mx0;
      buf_acc_data_5_4_0_sva <= buf_acc_data_5_4_0_sva_mx0;
      buf_acc_data_5_4_45_1_sva <= buf_acc_data_5_4_45_1_sva_mx0;
      buf_acc_data_5_4_56_46_sva <= buf_acc_data_5_4_56_46_sva_mx0;
      buf_acc_data_12_12_0_sva <= buf_acc_data_12_12_0_sva_mx0;
      buf_acc_data_12_12_45_1_sva <= buf_acc_data_12_12_45_1_sva_mx0;
      buf_acc_data_12_12_56_46_sva <= buf_acc_data_12_12_56_46_sva_mx0;
      buf_acc_data_5_5_0_sva <= buf_acc_data_5_5_0_sva_mx0;
      buf_acc_data_5_5_45_1_sva <= buf_acc_data_5_5_45_1_sva_mx0;
      buf_acc_data_5_5_56_46_sva <= buf_acc_data_5_5_56_46_sva_mx0;
      buf_acc_data_12_11_0_sva <= buf_acc_data_12_11_0_sva_mx0;
      buf_acc_data_12_11_45_1_sva <= buf_acc_data_12_11_45_1_sva_mx0;
      buf_acc_data_12_11_56_46_sva <= buf_acc_data_12_11_56_46_sva_mx0;
      buf_acc_data_5_6_0_sva <= buf_acc_data_5_6_0_sva_mx0;
      buf_acc_data_5_6_45_1_sva <= buf_acc_data_5_6_45_1_sva_mx0;
      buf_acc_data_5_6_56_46_sva <= buf_acc_data_5_6_56_46_sva_mx0;
      buf_acc_data_12_10_0_sva <= buf_acc_data_12_10_0_sva_mx0;
      buf_acc_data_12_10_45_1_sva <= buf_acc_data_12_10_45_1_sva_mx0;
      buf_acc_data_12_10_56_46_sva <= buf_acc_data_12_10_56_46_sva_mx0;
      buf_acc_data_5_7_0_sva <= buf_acc_data_5_7_0_sva_mx0;
      buf_acc_data_5_7_45_1_sva <= buf_acc_data_5_7_45_1_sva_mx0;
      buf_acc_data_5_7_56_46_sva <= buf_acc_data_5_7_56_46_sva_mx0;
      buf_acc_data_12_9_0_sva <= buf_acc_data_12_9_0_sva_mx0;
      buf_acc_data_12_9_45_1_sva <= buf_acc_data_12_9_45_1_sva_mx0;
      buf_acc_data_12_9_56_46_sva <= buf_acc_data_12_9_56_46_sva_mx0;
      buf_acc_data_5_8_0_sva <= buf_acc_data_5_8_0_sva_mx0;
      buf_acc_data_5_8_45_1_sva <= buf_acc_data_5_8_45_1_sva_mx0;
      buf_acc_data_5_8_56_46_sva <= buf_acc_data_5_8_56_46_sva_mx0;
      buf_acc_data_12_8_0_sva <= buf_acc_data_12_8_0_sva_mx0;
      buf_acc_data_12_8_45_1_sva <= buf_acc_data_12_8_45_1_sva_mx0;
      buf_acc_data_12_8_56_46_sva <= buf_acc_data_12_8_56_46_sva_mx0;
      buf_acc_data_5_9_0_sva <= buf_acc_data_5_9_0_sva_mx0;
      buf_acc_data_5_9_45_1_sva <= buf_acc_data_5_9_45_1_sva_mx0;
      buf_acc_data_5_9_56_46_sva <= buf_acc_data_5_9_56_46_sva_mx0;
      buf_acc_data_12_7_0_sva <= buf_acc_data_12_7_0_sva_mx0;
      buf_acc_data_12_7_45_1_sva <= buf_acc_data_12_7_45_1_sva_mx0;
      buf_acc_data_12_7_56_46_sva <= buf_acc_data_12_7_56_46_sva_mx0;
      buf_acc_data_5_10_0_sva <= buf_acc_data_5_10_0_sva_mx0;
      buf_acc_data_5_10_45_1_sva <= buf_acc_data_5_10_45_1_sva_mx0;
      buf_acc_data_5_10_56_46_sva <= buf_acc_data_5_10_56_46_sva_mx0;
      buf_acc_data_12_6_0_sva <= buf_acc_data_12_6_0_sva_mx0;
      buf_acc_data_12_6_45_1_sva <= buf_acc_data_12_6_45_1_sva_mx0;
      buf_acc_data_12_6_56_46_sva <= buf_acc_data_12_6_56_46_sva_mx0;
      buf_acc_data_5_11_0_sva <= buf_acc_data_5_11_0_sva_mx0;
      buf_acc_data_5_11_45_1_sva <= buf_acc_data_5_11_45_1_sva_mx0;
      buf_acc_data_5_11_56_46_sva <= buf_acc_data_5_11_56_46_sva_mx0;
      buf_acc_data_12_5_0_sva <= buf_acc_data_12_5_0_sva_mx0;
      buf_acc_data_12_5_45_1_sva <= buf_acc_data_12_5_45_1_sva_mx0;
      buf_acc_data_12_5_56_46_sva <= buf_acc_data_12_5_56_46_sva_mx0;
      buf_acc_data_5_12_0_sva <= buf_acc_data_5_12_0_sva_mx0;
      buf_acc_data_5_12_45_1_sva <= buf_acc_data_5_12_45_1_sva_mx0;
      buf_acc_data_5_12_56_46_sva <= buf_acc_data_5_12_56_46_sva_mx0;
      buf_acc_data_12_4_0_sva <= buf_acc_data_12_4_0_sva_mx0;
      buf_acc_data_12_4_45_1_sva <= buf_acc_data_12_4_45_1_sva_mx0;
      buf_acc_data_12_4_56_46_sva <= buf_acc_data_12_4_56_46_sva_mx0;
      buf_acc_data_5_13_0_sva <= buf_acc_data_5_13_0_sva_mx0;
      buf_acc_data_5_13_45_1_sva <= buf_acc_data_5_13_45_1_sva_mx0;
      buf_acc_data_5_13_56_46_sva <= buf_acc_data_5_13_56_46_sva_mx0;
      buf_acc_data_12_3_0_sva <= buf_acc_data_12_3_0_sva_mx0;
      buf_acc_data_12_3_45_1_sva <= buf_acc_data_12_3_45_1_sva_mx0;
      buf_acc_data_12_3_56_46_sva <= buf_acc_data_12_3_56_46_sva_mx0;
      buf_acc_data_5_14_0_sva <= buf_acc_data_5_14_0_sva_mx0;
      buf_acc_data_5_14_45_1_sva <= buf_acc_data_5_14_45_1_sva_mx0;
      buf_acc_data_5_14_56_46_sva <= buf_acc_data_5_14_56_46_sva_mx0;
      buf_acc_data_12_2_0_sva <= buf_acc_data_12_2_0_sva_mx0;
      buf_acc_data_12_2_45_1_sva <= buf_acc_data_12_2_45_1_sva_mx0;
      buf_acc_data_12_2_56_46_sva <= buf_acc_data_12_2_56_46_sva_mx0;
      buf_acc_data_5_15_0_sva <= buf_acc_data_5_15_0_sva_mx0;
      buf_acc_data_5_15_45_1_sva <= buf_acc_data_5_15_45_1_sva_mx0;
      buf_acc_data_5_15_56_46_sva <= buf_acc_data_5_15_56_46_sva_mx0;
      buf_acc_data_12_1_0_sva <= buf_acc_data_12_1_0_sva_mx0;
      buf_acc_data_12_1_45_1_sva <= buf_acc_data_12_1_45_1_sva_mx0;
      buf_acc_data_12_1_56_46_sva <= buf_acc_data_12_1_56_46_sva_mx0;
      buf_acc_data_5_16_0_sva <= buf_acc_data_5_16_0_sva_mx0;
      buf_acc_data_5_16_45_1_sva <= buf_acc_data_5_16_45_1_sva_mx0;
      buf_acc_data_5_16_56_46_sva <= buf_acc_data_5_16_56_46_sva_mx0;
      buf_acc_data_12_0_0_sva <= buf_acc_data_12_0_0_sva_mx0;
      buf_acc_data_12_0_45_1_sva <= buf_acc_data_12_0_45_1_sva_mx0;
      buf_acc_data_12_0_56_46_sva <= buf_acc_data_12_0_56_46_sva_mx0;
      buf_acc_data_5_17_0_sva <= buf_acc_data_5_17_0_sva_mx0;
      buf_acc_data_5_17_45_1_sva <= buf_acc_data_5_17_45_1_sva_mx0;
      buf_acc_data_5_17_56_46_sva <= buf_acc_data_5_17_56_46_sva_mx0;
      buf_acc_data_11_17_0_sva <= buf_acc_data_11_17_0_sva_mx0;
      buf_acc_data_11_17_45_1_sva <= buf_acc_data_11_17_45_1_sva_mx0;
      buf_acc_data_11_17_56_46_sva <= buf_acc_data_11_17_56_46_sva_mx0;
      buf_acc_data_6_0_0_sva <= buf_acc_data_6_0_0_sva_mx0;
      buf_acc_data_6_0_45_1_sva <= buf_acc_data_6_0_45_1_sva_mx0;
      buf_acc_data_6_0_56_46_sva <= buf_acc_data_6_0_56_46_sva_mx0;
      buf_acc_data_11_16_0_sva <= buf_acc_data_11_16_0_sva_mx0;
      buf_acc_data_11_16_45_1_sva <= buf_acc_data_11_16_45_1_sva_mx0;
      buf_acc_data_11_16_56_46_sva <= buf_acc_data_11_16_56_46_sva_mx0;
      buf_acc_data_6_1_0_sva <= buf_acc_data_6_1_0_sva_mx0;
      buf_acc_data_6_1_45_1_sva <= buf_acc_data_6_1_45_1_sva_mx0;
      buf_acc_data_6_1_56_46_sva <= buf_acc_data_6_1_56_46_sva_mx0;
      buf_acc_data_11_15_0_sva <= buf_acc_data_11_15_0_sva_mx0;
      buf_acc_data_11_15_45_1_sva <= buf_acc_data_11_15_45_1_sva_mx0;
      buf_acc_data_11_15_56_46_sva <= buf_acc_data_11_15_56_46_sva_mx0;
      buf_acc_data_6_2_0_sva <= buf_acc_data_6_2_0_sva_mx0;
      buf_acc_data_6_2_45_1_sva <= buf_acc_data_6_2_45_1_sva_mx0;
      buf_acc_data_6_2_56_46_sva <= buf_acc_data_6_2_56_46_sva_mx0;
      buf_acc_data_11_14_0_sva <= buf_acc_data_11_14_0_sva_mx0;
      buf_acc_data_11_14_45_1_sva <= buf_acc_data_11_14_45_1_sva_mx0;
      buf_acc_data_11_14_56_46_sva <= buf_acc_data_11_14_56_46_sva_mx0;
      buf_acc_data_6_3_0_sva <= buf_acc_data_6_3_0_sva_mx0;
      buf_acc_data_6_3_45_1_sva <= buf_acc_data_6_3_45_1_sva_mx0;
      buf_acc_data_6_3_56_46_sva <= buf_acc_data_6_3_56_46_sva_mx0;
      buf_acc_data_11_13_0_sva <= buf_acc_data_11_13_0_sva_mx0;
      buf_acc_data_11_13_45_1_sva <= buf_acc_data_11_13_45_1_sva_mx0;
      buf_acc_data_11_13_56_46_sva <= buf_acc_data_11_13_56_46_sva_mx0;
      buf_acc_data_6_4_0_sva <= buf_acc_data_6_4_0_sva_mx0;
      buf_acc_data_6_4_45_1_sva <= buf_acc_data_6_4_45_1_sva_mx0;
      buf_acc_data_6_4_56_46_sva <= buf_acc_data_6_4_56_46_sva_mx0;
      buf_acc_data_11_12_0_sva <= buf_acc_data_11_12_0_sva_mx0;
      buf_acc_data_11_12_45_1_sva <= buf_acc_data_11_12_45_1_sva_mx0;
      buf_acc_data_11_12_56_46_sva <= buf_acc_data_11_12_56_46_sva_mx0;
      buf_acc_data_6_5_0_sva <= buf_acc_data_6_5_0_sva_mx0;
      buf_acc_data_6_5_45_1_sva <= buf_acc_data_6_5_45_1_sva_mx0;
      buf_acc_data_6_5_56_46_sva <= buf_acc_data_6_5_56_46_sva_mx0;
      buf_acc_data_11_11_0_sva <= buf_acc_data_11_11_0_sva_mx0;
      buf_acc_data_11_11_45_1_sva <= buf_acc_data_11_11_45_1_sva_mx0;
      buf_acc_data_11_11_56_46_sva <= buf_acc_data_11_11_56_46_sva_mx0;
      buf_acc_data_6_6_0_sva <= buf_acc_data_6_6_0_sva_mx0;
      buf_acc_data_6_6_45_1_sva <= buf_acc_data_6_6_45_1_sva_mx0;
      buf_acc_data_6_6_56_46_sva <= buf_acc_data_6_6_56_46_sva_mx0;
      buf_acc_data_11_10_0_sva <= buf_acc_data_11_10_0_sva_mx0;
      buf_acc_data_11_10_45_1_sva <= buf_acc_data_11_10_45_1_sva_mx0;
      buf_acc_data_11_10_56_46_sva <= buf_acc_data_11_10_56_46_sva_mx0;
      buf_acc_data_6_7_0_sva <= buf_acc_data_6_7_0_sva_mx0;
      buf_acc_data_6_7_45_1_sva <= buf_acc_data_6_7_45_1_sva_mx0;
      buf_acc_data_6_7_56_46_sva <= buf_acc_data_6_7_56_46_sva_mx0;
      buf_acc_data_11_9_0_sva <= buf_acc_data_11_9_0_sva_mx0;
      buf_acc_data_11_9_45_1_sva <= buf_acc_data_11_9_45_1_sva_mx0;
      buf_acc_data_11_9_56_46_sva <= buf_acc_data_11_9_56_46_sva_mx0;
      buf_acc_data_6_8_0_sva <= buf_acc_data_6_8_0_sva_mx0;
      buf_acc_data_6_8_45_1_sva <= buf_acc_data_6_8_45_1_sva_mx0;
      buf_acc_data_6_8_56_46_sva <= buf_acc_data_6_8_56_46_sva_mx0;
      buf_acc_data_11_8_0_sva <= buf_acc_data_11_8_0_sva_mx0;
      buf_acc_data_11_8_45_1_sva <= buf_acc_data_11_8_45_1_sva_mx0;
      buf_acc_data_11_8_56_46_sva <= buf_acc_data_11_8_56_46_sva_mx0;
      buf_acc_data_6_9_0_sva <= buf_acc_data_6_9_0_sva_mx0;
      buf_acc_data_6_9_45_1_sva <= buf_acc_data_6_9_45_1_sva_mx0;
      buf_acc_data_6_9_56_46_sva <= buf_acc_data_6_9_56_46_sva_mx0;
      buf_acc_data_11_7_0_sva <= buf_acc_data_11_7_0_sva_mx0;
      buf_acc_data_11_7_45_1_sva <= buf_acc_data_11_7_45_1_sva_mx0;
      buf_acc_data_11_7_56_46_sva <= buf_acc_data_11_7_56_46_sva_mx0;
      buf_acc_data_6_10_0_sva <= buf_acc_data_6_10_0_sva_mx0;
      buf_acc_data_6_10_45_1_sva <= buf_acc_data_6_10_45_1_sva_mx0;
      buf_acc_data_6_10_56_46_sva <= buf_acc_data_6_10_56_46_sva_mx0;
      buf_acc_data_11_6_0_sva <= buf_acc_data_11_6_0_sva_mx0;
      buf_acc_data_11_6_45_1_sva <= buf_acc_data_11_6_45_1_sva_mx0;
      buf_acc_data_11_6_56_46_sva <= buf_acc_data_11_6_56_46_sva_mx0;
      buf_acc_data_6_11_0_sva <= buf_acc_data_6_11_0_sva_mx0;
      buf_acc_data_6_11_45_1_sva <= buf_acc_data_6_11_45_1_sva_mx0;
      buf_acc_data_6_11_56_46_sva <= buf_acc_data_6_11_56_46_sva_mx0;
      buf_acc_data_11_5_0_sva <= buf_acc_data_11_5_0_sva_mx0;
      buf_acc_data_11_5_45_1_sva <= buf_acc_data_11_5_45_1_sva_mx0;
      buf_acc_data_11_5_56_46_sva <= buf_acc_data_11_5_56_46_sva_mx0;
      buf_acc_data_6_12_0_sva <= buf_acc_data_6_12_0_sva_mx0;
      buf_acc_data_6_12_45_1_sva <= buf_acc_data_6_12_45_1_sva_mx0;
      buf_acc_data_6_12_56_46_sva <= buf_acc_data_6_12_56_46_sva_mx0;
      buf_acc_data_11_4_0_sva <= buf_acc_data_11_4_0_sva_mx0;
      buf_acc_data_11_4_45_1_sva <= buf_acc_data_11_4_45_1_sva_mx0;
      buf_acc_data_11_4_56_46_sva <= buf_acc_data_11_4_56_46_sva_mx0;
      buf_acc_data_6_13_0_sva <= buf_acc_data_6_13_0_sva_mx0;
      buf_acc_data_6_13_45_1_sva <= buf_acc_data_6_13_45_1_sva_mx0;
      buf_acc_data_6_13_56_46_sva <= buf_acc_data_6_13_56_46_sva_mx0;
      buf_acc_data_11_3_0_sva <= buf_acc_data_11_3_0_sva_mx0;
      buf_acc_data_11_3_45_1_sva <= buf_acc_data_11_3_45_1_sva_mx0;
      buf_acc_data_11_3_56_46_sva <= buf_acc_data_11_3_56_46_sva_mx0;
      buf_acc_data_6_14_0_sva <= buf_acc_data_6_14_0_sva_mx0;
      buf_acc_data_6_14_45_1_sva <= buf_acc_data_6_14_45_1_sva_mx0;
      buf_acc_data_6_14_56_46_sva <= buf_acc_data_6_14_56_46_sva_mx0;
      buf_acc_data_11_2_0_sva <= buf_acc_data_11_2_0_sva_mx0;
      buf_acc_data_11_2_45_1_sva <= buf_acc_data_11_2_45_1_sva_mx0;
      buf_acc_data_11_2_56_46_sva <= buf_acc_data_11_2_56_46_sva_mx0;
      buf_acc_data_6_15_0_sva <= buf_acc_data_6_15_0_sva_mx0;
      buf_acc_data_6_15_45_1_sva <= buf_acc_data_6_15_45_1_sva_mx0;
      buf_acc_data_6_15_56_46_sva <= buf_acc_data_6_15_56_46_sva_mx0;
      buf_acc_data_11_1_0_sva <= buf_acc_data_11_1_0_sva_mx0;
      buf_acc_data_11_1_45_1_sva <= buf_acc_data_11_1_45_1_sva_mx0;
      buf_acc_data_11_1_56_46_sva <= buf_acc_data_11_1_56_46_sva_mx0;
      buf_acc_data_6_16_0_sva <= buf_acc_data_6_16_0_sva_mx0;
      buf_acc_data_6_16_45_1_sva <= buf_acc_data_6_16_45_1_sva_mx0;
      buf_acc_data_6_16_56_46_sva <= buf_acc_data_6_16_56_46_sva_mx0;
      buf_acc_data_11_0_0_sva <= buf_acc_data_11_0_0_sva_mx0;
      buf_acc_data_11_0_45_1_sva <= buf_acc_data_11_0_45_1_sva_mx0;
      buf_acc_data_11_0_56_46_sva <= buf_acc_data_11_0_56_46_sva_mx0;
      buf_acc_data_6_17_0_sva <= buf_acc_data_6_17_0_sva_mx0;
      buf_acc_data_6_17_45_1_sva <= buf_acc_data_6_17_45_1_sva_mx0;
      buf_acc_data_6_17_56_46_sva <= buf_acc_data_6_17_56_46_sva_mx0;
      buf_acc_data_10_17_0_sva <= buf_acc_data_10_17_0_sva_mx0;
      buf_acc_data_10_17_45_1_sva <= buf_acc_data_10_17_45_1_sva_mx0;
      buf_acc_data_10_17_56_46_sva <= buf_acc_data_10_17_56_46_sva_mx0;
      buf_acc_data_7_0_0_sva <= buf_acc_data_7_0_0_sva_mx0;
      buf_acc_data_7_0_45_1_sva <= buf_acc_data_7_0_45_1_sva_mx0;
      buf_acc_data_7_0_56_46_sva <= buf_acc_data_7_0_56_46_sva_mx0;
      buf_acc_data_10_16_0_sva <= buf_acc_data_10_16_0_sva_mx0;
      buf_acc_data_10_16_45_1_sva <= buf_acc_data_10_16_45_1_sva_mx0;
      buf_acc_data_10_16_56_46_sva <= buf_acc_data_10_16_56_46_sva_mx0;
      buf_acc_data_7_1_0_sva <= buf_acc_data_7_1_0_sva_mx0;
      buf_acc_data_7_1_45_1_sva <= buf_acc_data_7_1_45_1_sva_mx0;
      buf_acc_data_7_1_56_46_sva <= buf_acc_data_7_1_56_46_sva_mx0;
      buf_acc_data_10_15_0_sva <= buf_acc_data_10_15_0_sva_mx0;
      buf_acc_data_10_15_45_1_sva <= buf_acc_data_10_15_45_1_sva_mx0;
      buf_acc_data_10_15_56_46_sva <= buf_acc_data_10_15_56_46_sva_mx0;
      buf_acc_data_7_2_0_sva <= buf_acc_data_7_2_0_sva_mx0;
      buf_acc_data_7_2_45_1_sva <= buf_acc_data_7_2_45_1_sva_mx0;
      buf_acc_data_7_2_56_46_sva <= buf_acc_data_7_2_56_46_sva_mx0;
      buf_acc_data_10_14_0_sva <= buf_acc_data_10_14_0_sva_mx0;
      buf_acc_data_10_14_45_1_sva <= buf_acc_data_10_14_45_1_sva_mx0;
      buf_acc_data_10_14_56_46_sva <= buf_acc_data_10_14_56_46_sva_mx0;
      buf_acc_data_7_3_0_sva <= buf_acc_data_7_3_0_sva_mx0;
      buf_acc_data_7_3_45_1_sva <= buf_acc_data_7_3_45_1_sva_mx0;
      buf_acc_data_7_3_56_46_sva <= buf_acc_data_7_3_56_46_sva_mx0;
      buf_acc_data_10_13_0_sva <= buf_acc_data_10_13_0_sva_mx0;
      buf_acc_data_10_13_45_1_sva <= buf_acc_data_10_13_45_1_sva_mx0;
      buf_acc_data_10_13_56_46_sva <= buf_acc_data_10_13_56_46_sva_mx0;
      buf_acc_data_7_4_0_sva <= buf_acc_data_7_4_0_sva_mx0;
      buf_acc_data_7_4_45_1_sva <= buf_acc_data_7_4_45_1_sva_mx0;
      buf_acc_data_7_4_56_46_sva <= buf_acc_data_7_4_56_46_sva_mx0;
      buf_acc_data_10_12_0_sva <= buf_acc_data_10_12_0_sva_mx0;
      buf_acc_data_10_12_45_1_sva <= buf_acc_data_10_12_45_1_sva_mx0;
      buf_acc_data_10_12_56_46_sva <= buf_acc_data_10_12_56_46_sva_mx0;
      buf_acc_data_7_5_0_sva <= buf_acc_data_7_5_0_sva_mx0;
      buf_acc_data_7_5_45_1_sva <= buf_acc_data_7_5_45_1_sva_mx0;
      buf_acc_data_7_5_56_46_sva <= buf_acc_data_7_5_56_46_sva_mx0;
      buf_acc_data_10_11_0_sva <= buf_acc_data_10_11_0_sva_mx0;
      buf_acc_data_10_11_45_1_sva <= buf_acc_data_10_11_45_1_sva_mx0;
      buf_acc_data_10_11_56_46_sva <= buf_acc_data_10_11_56_46_sva_mx0;
      buf_acc_data_7_6_0_sva <= buf_acc_data_7_6_0_sva_mx0;
      buf_acc_data_7_6_45_1_sva <= buf_acc_data_7_6_45_1_sva_mx0;
      buf_acc_data_7_6_56_46_sva <= buf_acc_data_7_6_56_46_sva_mx0;
      buf_acc_data_10_10_0_sva <= buf_acc_data_10_10_0_sva_mx0;
      buf_acc_data_10_10_45_1_sva <= buf_acc_data_10_10_45_1_sva_mx0;
      buf_acc_data_10_10_56_46_sva <= buf_acc_data_10_10_56_46_sva_mx0;
      buf_acc_data_7_7_0_sva <= buf_acc_data_7_7_0_sva_mx0;
      buf_acc_data_7_7_45_1_sva <= buf_acc_data_7_7_45_1_sva_mx0;
      buf_acc_data_7_7_56_46_sva <= buf_acc_data_7_7_56_46_sva_mx0;
      buf_acc_data_10_9_0_sva <= buf_acc_data_10_9_0_sva_mx0;
      buf_acc_data_10_9_45_1_sva <= buf_acc_data_10_9_45_1_sva_mx0;
      buf_acc_data_10_9_56_46_sva <= buf_acc_data_10_9_56_46_sva_mx0;
      buf_acc_data_7_8_0_sva <= buf_acc_data_7_8_0_sva_mx0;
      buf_acc_data_7_8_45_1_sva <= buf_acc_data_7_8_45_1_sva_mx0;
      buf_acc_data_7_8_56_46_sva <= buf_acc_data_7_8_56_46_sva_mx0;
      buf_acc_data_10_8_0_sva <= buf_acc_data_10_8_0_sva_mx0;
      buf_acc_data_10_8_45_1_sva <= buf_acc_data_10_8_45_1_sva_mx0;
      buf_acc_data_10_8_56_46_sva <= buf_acc_data_10_8_56_46_sva_mx0;
      buf_acc_data_7_9_0_sva <= buf_acc_data_7_9_0_sva_mx0;
      buf_acc_data_7_9_45_1_sva <= buf_acc_data_7_9_45_1_sva_mx0;
      buf_acc_data_7_9_56_46_sva <= buf_acc_data_7_9_56_46_sva_mx0;
      buf_acc_data_10_7_0_sva <= buf_acc_data_10_7_0_sva_mx0;
      buf_acc_data_10_7_45_1_sva <= buf_acc_data_10_7_45_1_sva_mx0;
      buf_acc_data_10_7_56_46_sva <= buf_acc_data_10_7_56_46_sva_mx0;
      buf_acc_data_7_10_0_sva <= buf_acc_data_7_10_0_sva_mx0;
      buf_acc_data_7_10_45_1_sva <= buf_acc_data_7_10_45_1_sva_mx0;
      buf_acc_data_7_10_56_46_sva <= buf_acc_data_7_10_56_46_sva_mx0;
      buf_acc_data_10_6_0_sva <= buf_acc_data_10_6_0_sva_mx0;
      buf_acc_data_10_6_45_1_sva <= buf_acc_data_10_6_45_1_sva_mx0;
      buf_acc_data_10_6_56_46_sva <= buf_acc_data_10_6_56_46_sva_mx0;
      buf_acc_data_7_11_0_sva <= buf_acc_data_7_11_0_sva_mx0;
      buf_acc_data_7_11_45_1_sva <= buf_acc_data_7_11_45_1_sva_mx0;
      buf_acc_data_7_11_56_46_sva <= buf_acc_data_7_11_56_46_sva_mx0;
      buf_acc_data_10_5_0_sva <= buf_acc_data_10_5_0_sva_mx0;
      buf_acc_data_10_5_45_1_sva <= buf_acc_data_10_5_45_1_sva_mx0;
      buf_acc_data_10_5_56_46_sva <= buf_acc_data_10_5_56_46_sva_mx0;
      buf_acc_data_7_12_0_sva <= buf_acc_data_7_12_0_sva_mx0;
      buf_acc_data_7_12_45_1_sva <= buf_acc_data_7_12_45_1_sva_mx0;
      buf_acc_data_7_12_56_46_sva <= buf_acc_data_7_12_56_46_sva_mx0;
      buf_acc_data_10_4_0_sva <= buf_acc_data_10_4_0_sva_mx0;
      buf_acc_data_10_4_45_1_sva <= buf_acc_data_10_4_45_1_sva_mx0;
      buf_acc_data_10_4_56_46_sva <= buf_acc_data_10_4_56_46_sva_mx0;
      buf_acc_data_7_13_0_sva <= buf_acc_data_7_13_0_sva_mx0;
      buf_acc_data_7_13_45_1_sva <= buf_acc_data_7_13_45_1_sva_mx0;
      buf_acc_data_7_13_56_46_sva <= buf_acc_data_7_13_56_46_sva_mx0;
      buf_acc_data_10_3_0_sva <= buf_acc_data_10_3_0_sva_mx0;
      buf_acc_data_10_3_45_1_sva <= buf_acc_data_10_3_45_1_sva_mx0;
      buf_acc_data_10_3_56_46_sva <= buf_acc_data_10_3_56_46_sva_mx0;
      buf_acc_data_7_14_0_sva <= buf_acc_data_7_14_0_sva_mx0;
      buf_acc_data_7_14_45_1_sva <= buf_acc_data_7_14_45_1_sva_mx0;
      buf_acc_data_7_14_56_46_sva <= buf_acc_data_7_14_56_46_sva_mx0;
      buf_acc_data_10_2_0_sva <= buf_acc_data_10_2_0_sva_mx0;
      buf_acc_data_10_2_45_1_sva <= buf_acc_data_10_2_45_1_sva_mx0;
      buf_acc_data_10_2_56_46_sva <= buf_acc_data_10_2_56_46_sva_mx0;
      buf_acc_data_7_15_0_sva <= buf_acc_data_7_15_0_sva_mx0;
      buf_acc_data_7_15_45_1_sva <= buf_acc_data_7_15_45_1_sva_mx0;
      buf_acc_data_7_15_56_46_sva <= buf_acc_data_7_15_56_46_sva_mx0;
      buf_acc_data_10_1_0_sva <= buf_acc_data_10_1_0_sva_mx0;
      buf_acc_data_10_1_45_1_sva <= buf_acc_data_10_1_45_1_sva_mx0;
      buf_acc_data_10_1_56_46_sva <= buf_acc_data_10_1_56_46_sva_mx0;
      buf_acc_data_7_16_0_sva <= buf_acc_data_7_16_0_sva_mx0;
      buf_acc_data_7_16_45_1_sva <= buf_acc_data_7_16_45_1_sva_mx0;
      buf_acc_data_7_16_56_46_sva <= buf_acc_data_7_16_56_46_sva_mx0;
      buf_acc_data_10_0_0_sva <= buf_acc_data_10_0_0_sva_mx0;
      buf_acc_data_10_0_45_1_sva <= buf_acc_data_10_0_45_1_sva_mx0;
      buf_acc_data_10_0_56_46_sva <= buf_acc_data_10_0_56_46_sva_mx0;
      buf_acc_data_7_17_0_sva <= buf_acc_data_7_17_0_sva_mx0;
      buf_acc_data_7_17_45_1_sva <= buf_acc_data_7_17_45_1_sva_mx0;
      buf_acc_data_7_17_56_46_sva <= buf_acc_data_7_17_56_46_sva_mx0;
      buf_acc_data_9_17_0_sva <= buf_acc_data_9_17_0_sva_mx0;
      buf_acc_data_9_17_45_1_sva <= buf_acc_data_9_17_45_1_sva_mx0;
      buf_acc_data_9_17_56_46_sva <= buf_acc_data_9_17_56_46_sva_mx0;
      buf_acc_data_8_0_0_sva <= buf_acc_data_8_0_0_sva_mx0;
      buf_acc_data_8_0_45_1_sva <= buf_acc_data_8_0_45_1_sva_mx0;
      buf_acc_data_8_0_56_46_sva <= buf_acc_data_8_0_56_46_sva_mx0;
      buf_acc_data_9_16_0_sva <= buf_acc_data_9_16_0_sva_mx0;
      buf_acc_data_9_16_45_1_sva <= buf_acc_data_9_16_45_1_sva_mx0;
      buf_acc_data_9_16_56_46_sva <= buf_acc_data_9_16_56_46_sva_mx0;
      buf_acc_data_8_1_0_sva <= buf_acc_data_8_1_0_sva_mx0;
      buf_acc_data_8_1_45_1_sva <= buf_acc_data_8_1_45_1_sva_mx0;
      buf_acc_data_8_1_56_46_sva <= buf_acc_data_8_1_56_46_sva_mx0;
      buf_acc_data_9_15_0_sva <= buf_acc_data_9_15_0_sva_mx0;
      buf_acc_data_9_15_45_1_sva <= buf_acc_data_9_15_45_1_sva_mx0;
      buf_acc_data_9_15_56_46_sva <= buf_acc_data_9_15_56_46_sva_mx0;
      buf_acc_data_8_2_0_sva <= buf_acc_data_8_2_0_sva_mx0;
      buf_acc_data_8_2_45_1_sva <= buf_acc_data_8_2_45_1_sva_mx0;
      buf_acc_data_8_2_56_46_sva <= buf_acc_data_8_2_56_46_sva_mx0;
      buf_acc_data_9_14_0_sva <= buf_acc_data_9_14_0_sva_mx0;
      buf_acc_data_9_14_45_1_sva <= buf_acc_data_9_14_45_1_sva_mx0;
      buf_acc_data_9_14_56_46_sva <= buf_acc_data_9_14_56_46_sva_mx0;
      buf_acc_data_8_3_0_sva <= buf_acc_data_8_3_0_sva_mx0;
      buf_acc_data_8_3_45_1_sva <= buf_acc_data_8_3_45_1_sva_mx0;
      buf_acc_data_8_3_56_46_sva <= buf_acc_data_8_3_56_46_sva_mx0;
      buf_acc_data_9_13_0_sva <= buf_acc_data_9_13_0_sva_mx0;
      buf_acc_data_9_13_45_1_sva <= buf_acc_data_9_13_45_1_sva_mx0;
      buf_acc_data_9_13_56_46_sva <= buf_acc_data_9_13_56_46_sva_mx0;
      buf_acc_data_8_4_0_sva <= buf_acc_data_8_4_0_sva_mx0;
      buf_acc_data_8_4_45_1_sva <= buf_acc_data_8_4_45_1_sva_mx0;
      buf_acc_data_8_4_56_46_sva <= buf_acc_data_8_4_56_46_sva_mx0;
      buf_acc_data_9_12_0_sva <= buf_acc_data_9_12_0_sva_mx0;
      buf_acc_data_9_12_45_1_sva <= buf_acc_data_9_12_45_1_sva_mx0;
      buf_acc_data_9_12_56_46_sva <= buf_acc_data_9_12_56_46_sva_mx0;
      buf_acc_data_8_5_0_sva <= buf_acc_data_8_5_0_sva_mx0;
      buf_acc_data_8_5_45_1_sva <= buf_acc_data_8_5_45_1_sva_mx0;
      buf_acc_data_8_5_56_46_sva <= buf_acc_data_8_5_56_46_sva_mx0;
      buf_acc_data_9_11_0_sva <= buf_acc_data_9_11_0_sva_mx0;
      buf_acc_data_9_11_45_1_sva <= buf_acc_data_9_11_45_1_sva_mx0;
      buf_acc_data_9_11_56_46_sva <= buf_acc_data_9_11_56_46_sva_mx0;
      buf_acc_data_8_6_0_sva <= buf_acc_data_8_6_0_sva_mx0;
      buf_acc_data_8_6_45_1_sva <= buf_acc_data_8_6_45_1_sva_mx0;
      buf_acc_data_8_6_56_46_sva <= buf_acc_data_8_6_56_46_sva_mx0;
      buf_acc_data_9_10_0_sva <= buf_acc_data_9_10_0_sva_mx0;
      buf_acc_data_9_10_45_1_sva <= buf_acc_data_9_10_45_1_sva_mx0;
      buf_acc_data_9_10_56_46_sva <= buf_acc_data_9_10_56_46_sva_mx0;
      buf_acc_data_8_7_0_sva <= buf_acc_data_8_7_0_sva_mx0;
      buf_acc_data_8_7_45_1_sva <= buf_acc_data_8_7_45_1_sva_mx0;
      buf_acc_data_8_7_56_46_sva <= buf_acc_data_8_7_56_46_sva_mx0;
      buf_acc_data_9_9_0_sva <= buf_acc_data_9_9_0_sva_mx0;
      buf_acc_data_9_9_45_1_sva <= buf_acc_data_9_9_45_1_sva_mx0;
      buf_acc_data_9_9_56_46_sva <= buf_acc_data_9_9_56_46_sva_mx0;
      buf_acc_data_8_8_0_sva <= buf_acc_data_8_8_0_sva_mx0;
      buf_acc_data_8_8_45_1_sva <= buf_acc_data_8_8_45_1_sva_mx0;
      buf_acc_data_8_8_56_46_sva <= buf_acc_data_8_8_56_46_sva_mx0;
      buf_acc_data_9_8_0_sva <= buf_acc_data_9_8_0_sva_mx0;
      buf_acc_data_9_8_45_1_sva <= buf_acc_data_9_8_45_1_sva_mx0;
      buf_acc_data_9_8_56_46_sva <= buf_acc_data_9_8_56_46_sva_mx0;
      buf_acc_data_8_9_0_sva <= buf_acc_data_8_9_0_sva_mx0;
      buf_acc_data_8_9_45_1_sva <= buf_acc_data_8_9_45_1_sva_mx0;
      buf_acc_data_8_9_56_46_sva <= buf_acc_data_8_9_56_46_sva_mx0;
      buf_acc_data_9_7_0_sva <= buf_acc_data_9_7_0_sva_mx0;
      buf_acc_data_9_7_45_1_sva <= buf_acc_data_9_7_45_1_sva_mx0;
      buf_acc_data_9_7_56_46_sva <= buf_acc_data_9_7_56_46_sva_mx0;
      buf_acc_data_8_10_0_sva <= buf_acc_data_8_10_0_sva_mx0;
      buf_acc_data_8_10_45_1_sva <= buf_acc_data_8_10_45_1_sva_mx0;
      buf_acc_data_8_10_56_46_sva <= buf_acc_data_8_10_56_46_sva_mx0;
      buf_acc_data_9_6_0_sva <= buf_acc_data_9_6_0_sva_mx0;
      buf_acc_data_9_6_45_1_sva <= buf_acc_data_9_6_45_1_sva_mx0;
      buf_acc_data_9_6_56_46_sva <= buf_acc_data_9_6_56_46_sva_mx0;
      buf_acc_data_8_11_0_sva <= buf_acc_data_8_11_0_sva_mx0;
      buf_acc_data_8_11_45_1_sva <= buf_acc_data_8_11_45_1_sva_mx0;
      buf_acc_data_8_11_56_46_sva <= buf_acc_data_8_11_56_46_sva_mx0;
      buf_acc_data_9_5_0_sva <= buf_acc_data_9_5_0_sva_mx0;
      buf_acc_data_9_5_45_1_sva <= buf_acc_data_9_5_45_1_sva_mx0;
      buf_acc_data_9_5_56_46_sva <= buf_acc_data_9_5_56_46_sva_mx0;
      buf_acc_data_8_12_0_sva <= buf_acc_data_8_12_0_sva_mx0;
      buf_acc_data_8_12_45_1_sva <= buf_acc_data_8_12_45_1_sva_mx0;
      buf_acc_data_8_12_56_46_sva <= buf_acc_data_8_12_56_46_sva_mx0;
      buf_acc_data_9_4_0_sva <= buf_acc_data_9_4_0_sva_mx0;
      buf_acc_data_9_4_45_1_sva <= buf_acc_data_9_4_45_1_sva_mx0;
      buf_acc_data_9_4_56_46_sva <= buf_acc_data_9_4_56_46_sva_mx0;
      buf_acc_data_8_13_0_sva <= buf_acc_data_8_13_0_sva_mx0;
      buf_acc_data_8_13_45_1_sva <= buf_acc_data_8_13_45_1_sva_mx0;
      buf_acc_data_8_13_56_46_sva <= buf_acc_data_8_13_56_46_sva_mx0;
      buf_acc_data_9_3_0_sva <= buf_acc_data_9_3_0_sva_mx0;
      buf_acc_data_9_3_45_1_sva <= buf_acc_data_9_3_45_1_sva_mx0;
      buf_acc_data_9_3_56_46_sva <= buf_acc_data_9_3_56_46_sva_mx0;
      buf_acc_data_8_14_0_sva <= buf_acc_data_8_14_0_sva_mx0;
      buf_acc_data_8_14_45_1_sva <= buf_acc_data_8_14_45_1_sva_mx0;
      buf_acc_data_8_14_56_46_sva <= buf_acc_data_8_14_56_46_sva_mx0;
      buf_acc_data_9_2_0_sva <= buf_acc_data_9_2_0_sva_mx0;
      buf_acc_data_9_2_45_1_sva <= buf_acc_data_9_2_45_1_sva_mx0;
      buf_acc_data_9_2_56_46_sva <= buf_acc_data_9_2_56_46_sva_mx0;
      buf_acc_data_8_15_0_sva <= buf_acc_data_8_15_0_sva_mx0;
      buf_acc_data_8_15_45_1_sva <= buf_acc_data_8_15_45_1_sva_mx0;
      buf_acc_data_8_15_56_46_sva <= buf_acc_data_8_15_56_46_sva_mx0;
      buf_acc_data_9_1_0_sva <= buf_acc_data_9_1_0_sva_mx0;
      buf_acc_data_9_1_45_1_sva <= buf_acc_data_9_1_45_1_sva_mx0;
      buf_acc_data_9_1_56_46_sva <= buf_acc_data_9_1_56_46_sva_mx0;
      buf_acc_data_8_16_0_sva <= buf_acc_data_8_16_0_sva_mx0;
      buf_acc_data_8_16_45_1_sva <= buf_acc_data_8_16_45_1_sva_mx0;
      buf_acc_data_8_16_56_46_sva <= buf_acc_data_8_16_56_46_sva_mx0;
      buf_acc_data_9_0_0_sva <= buf_acc_data_9_0_0_sva_mx0;
      buf_acc_data_9_0_45_1_sva <= buf_acc_data_9_0_45_1_sva_mx0;
      buf_acc_data_9_0_56_46_sva <= buf_acc_data_9_0_56_46_sva_mx0;
      buf_acc_data_8_17_0_sva <= buf_acc_data_8_17_0_sva_mx0;
      buf_acc_data_8_17_45_1_sva <= buf_acc_data_8_17_45_1_sva_mx0;
      buf_acc_data_8_17_56_46_sva <= buf_acc_data_8_17_56_46_sva_mx0;
      CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2 <= MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_dfm_1,
          CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_mx1, fsm_output[2]);
      CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2 <= MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_dfm_1,
          CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_mx1, fsm_output[2]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_write_chnl_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_685 | or_tmp_676) ) begin
      reg_dma_write_chnl_rsci_ivld_core_psct_cse <= ~ or_tmp_685;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_read_chnl_rsci_irdy_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (((~ mux_331_nl) & BATCH_LOOP_and_6_tmp & (fsm_output[2]))
        | or_tmp_693) ) begin
      reg_dma_read_chnl_rsci_irdy_core_psct_cse <= ~ or_tmp_693;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_write_ctrl_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((or_316_cse & or_453_cse & nor_291_cse & BATCH_LOOP_and_6_tmp
        & (fsm_output[2])) | or_tmp_700) ) begin
      reg_dma_write_ctrl_rsci_ivld_core_psct_cse <= ~ or_tmp_700;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0 <= 1'b0;
      LOAD_LOOP_i_lpi_2_dfm_2 <= 16'b0000000000000000;
    end
    else if ( STORE_LOOP_and_703_cse ) begin
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2 <= reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1 <= reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0 <= reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse;
      LOAD_LOOP_i_lpi_2_dfm_2 <= LOAD_LOOP_i_lpi_2_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
          <= 1'b0;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_if_1_and_cse ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
          <= CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_2;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2 <= lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1 <= lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_1;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0 <= lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_2 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_1 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_0 <= 1'b0;
    end
    else if ( STORE_LOOP_and_709_cse ) begin
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_2 <= lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_1 <= lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1;
      lfst_exit_STORE_LOOP_lpi_2_dfm_st_4_0 <= lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_info_index_15_0_lpi_2 <= 16'b0000000000000000;
    end
    else if ( core_wen & ((mux_tmp_354 & BATCH_LOOP_and_6_tmp & (fsm_output[2]))
        | (fsm_output[3])) ) begin
      dma_read_info_index_15_0_lpi_2 <= MUX_v_16_2_2(z_out_6, dma_read_info_index_15_0_lpi_2_dfm,
          fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_chan_5_0_lpi_2_4_0 <= 5'b00000;
      CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0 <= 5'b00000;
    end
    else if ( PADDING_LOOP_chan_and_4_cse ) begin
      PADDING_LOOP_chan_5_0_lpi_2_4_0 <= MUX_v_5_2_2(PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0_mx1w0,
          PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0, fsm_output[3]);
      CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0 <= MUX_v_5_2_2(CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0_mx1w0,
          CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_PADDING_LOOP_for_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | mux_tmp_357 | (~ BATCH_LOOP_and_6_tmp)))
        ) begin
      exit_PADDING_LOOP_for_lpi_2_dfm_1 <= exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm <= 1'b0;
    end
    else if ( core_wen & (fsm_output[2]) & or_453_cse & nor_291_cse & BATCH_LOOP_and_6_tmp
        ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm <= exit_CONVOLUTION_LOOP_lpi_2_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | and_769_cse | and_770_cse | mux_325_cse
        | (~ BATCH_LOOP_and_6_tmp))) ) begin
      exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1 <= exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | and_770_cse | mux_325_cse | (~
        BATCH_LOOP_and_6_tmp))) ) begin
      exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1 <= exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | and_765_cse | mux_376_cse | (~
        BATCH_LOOP_and_6_tmp))) ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_STORE_LOOP_lpi_2_2 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_0 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2 <= 45'b000000000000000000000000000000000000000000000;
    end
    else if ( PADDING_LOOP_chan_and_cse ) begin
      lfst_exit_STORE_LOOP_lpi_2_2 <= MUX_s_1_2_2(lfst_exit_STORE_LOOP_lpi_2_2_mx1,
          lfst_exit_STORE_LOOP_lpi_2_dfm_8_2, fsm_output[3]);
      lfst_exit_STORE_LOOP_lpi_2_0 <= MUX_s_1_2_2(lfst_exit_STORE_LOOP_lpi_2_0_mx1,
          lfst_exit_STORE_LOOP_lpi_2_dfm_8_0, fsm_output[3]);
      lfst_exit_STORE_LOOP_lpi_2_1 <= MUX_s_1_2_2(lfst_exit_STORE_LOOP_lpi_2_1_mx1,
          lfst_exit_STORE_LOOP_lpi_2_dfm_8_1, fsm_output[3]);
      CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2 <= MUX_v_45_2_2(CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_mx1,
          CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_dfm_1, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_for_for_land_2_lpi_2_dfm_1 <= 1'b0;
      PADDING_LOOP_for_for_index_in_acc_itm_1 <= 14'b00000000000000;
      LOAD_LOOP_i_sva_1_1 <= 16'b0000000000000000;
    end
    else if ( PADDING_LOOP_for_for_aelse_2_and_2_cse ) begin
      PADDING_LOOP_for_for_land_2_lpi_2_dfm_1 <= PADDING_LOOP_for_for_land_2_lpi_2_dfm_mx1w0;
      PADDING_LOOP_for_for_index_in_acc_itm_1 <= nl_PADDING_LOOP_for_for_index_in_acc_itm_1[13:0];
      LOAD_LOOP_i_sva_1_1 <= z_out_12[15:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1 <= 1'b0;
    end
    else if ( core_wen & ((mux_378_nl & BATCH_LOOP_and_6_tmp & (fsm_output[2])) |
        PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1_mx0c1) ) begin
      PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1 <= MUX_s_1_2_2(PADDING_LOOP_for_for_land_2_lpi_2_dfm_mx1w0,
          PADDING_LOOP_for_for_land_2_lpi_2_dfm_st, PADDING_LOOP_for_for_land_2_lpi_2_dfm_st_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_k_slc_CONVOLUTION_LOOP_for_k_5_0_4_0_3_itm_1 <= 5'b00000;
    end
    else if ( core_wen & (((~(STORE_LOOP_or_2336_tmp | BATCH_LOOP_asn_itm_1)) & BATCH_LOOP_and_4_tmp
        & BATCH_LOOP_and_6_tmp & (fsm_output[2])) | and_148_rgt) ) begin
      CONVOLUTION_LOOP_for_k_slc_CONVOLUTION_LOOP_for_k_5_0_4_0_3_itm_1 <= MUX_v_5_2_2(CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0,
          CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0, and_148_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_760 | exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1_mx0c1)
        ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1 <= MUX_s_1_2_2(exit_CONVOLUTION_LOOP_lpi_2_dfm_2_mx0w0,
          exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st, exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_760 | exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1_mx0c1)
        ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1 <= MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1,
          exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st, exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1 <= 14'b00000000000000;
      CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1 <= 16'b0000000000000000;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_for_for_and_10_cse ) begin
      CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1 <= nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1[13:0];
      CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1 <= nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1[15:0];
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1 <= exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_BATCH_LOOP_lpi_2_dfm_2_1 <= 1'b0;
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0 <= 5'b00000;
    end
    else if ( BATCH_LOOP_and_14_cse ) begin
      exit_BATCH_LOOP_lpi_2_dfm_2_1 <= exit_BATCH_LOOP_lpi_2_dfm_2_mx1w0;
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_1_4_0 <= CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      BATCH_LOOP_asn_itm_1 <= 1'b0;
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse <= 1'b0;
      STORE_LOOP_and_35_itm_1 <= 1'b0;
      STORE_LOOP_or_tmp_1 <= 1'b0;
      STORE_LOOP_and_30_itm_1 <= 1'b0;
      STORE_LOOP_and_32_itm_1 <= 1'b0;
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse <= 1'b0;
      STORE_LOOP_or_2332_itm_1 <= 1'b0;
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse <= 1'b0;
      STORE_LOOP_equal_tmp_2_1 <= 1'b0;
      STORE_LOOP_and_15_itm_1 <= 1'b0;
      STORE_LOOP_or_2_itm_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_1_0 <= 1'b0;
      STORE_LOOP_data_asn_itm_1 <= 14'b00000000000000;
      PADDING_LOOP_for_row_4_0_lpi_2_dfm_5 <= 5'b00000;
      lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1 <= 1'b0;
      PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4 <= 5'b00000;
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0 <= 5'b00000;
      lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2 <= 8'b00000000;
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4 <= 3'b000;
      STORE_LOOP_i_13_0_lpi_2_dfm_2 <= 14'b00000000000000;
    end
    else if ( BATCH_LOOP_and_10_cse ) begin
      BATCH_LOOP_asn_itm_1 <= exit_BATCH_LOOP_lpi_2_dfm_2_mx1w0;
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_2_cse <= lfst_exit_STORE_LOOP_lpi_2_dfm_2_mx1w0;
      STORE_LOOP_and_35_itm_1 <= STORE_LOOP_and_tmp_1 & STORE_LOOP_equal_tmp_4;
      STORE_LOOP_or_tmp_1 <= STORE_LOOP_or_tmp_mx0w0;
      STORE_LOOP_and_30_itm_1 <= STORE_LOOP_and_30_cse;
      STORE_LOOP_and_32_itm_1 <= STORE_LOOP_and_32_cse;
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse <= lfst_exit_STORE_LOOP_lpi_2_dfm_0_mx0w1;
      STORE_LOOP_or_2332_itm_1 <= STORE_LOOP_and_29_cse | STORE_LOOP_and_31_cse |
          STORE_LOOP_and_33_cse | ((~ STORE_LOOP_and_tmp_1) & STORE_LOOP_equal_tmp_4)
          | STORE_LOOP_or_tmp_2;
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_1_cse <= lfst_exit_STORE_LOOP_lpi_2_dfm_1_mx0w1;
      STORE_LOOP_equal_tmp_2_1 <= STORE_LOOP_equal_tmp_2_mx0w0;
      STORE_LOOP_and_15_itm_1 <= (~ LOAD_LOOP_LOAD_LOOP_if_and_tmp) & STORE_LOOP_equal_tmp_6;
      STORE_LOOP_or_2_itm_1 <= (LOAD_LOOP_LOAD_LOOP_if_and_tmp & STORE_LOOP_equal_tmp_6)
          | STORE_LOOP_equal_tmp_5 | STORE_LOOP_equal_tmp_2_mx0w0 | STORE_LOOP_equal_tmp_4
          | STORE_LOOP_or_tmp_2;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_1_0 <= MUX_s_1_2_2((CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6[0]),
          reg_CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_ftd_4, mux_tmp_468);
      STORE_LOOP_data_asn_itm_1 <= STORE_LOOP_i_13_0_lpi_2;
      PADDING_LOOP_for_row_4_0_lpi_2_dfm_5 <= PADDING_LOOP_for_row_4_0_lpi_2_dfm_5_mx0w0;
      lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1 <= lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0;
      PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4 <= PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4_mx0w0;
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0 <= CONVOLUTION_LOOP_for_k_5_0_lpi_2_dfm_5_4_0_mx1w0;
      lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1 <= lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0;
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5 <= CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5_mx0w0;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5 <= CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5_mx0w0;
      CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2 <= CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2_mx0w0;
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3 <= CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3_mx0w0;
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4 <= CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4_mx0w0;
      STORE_LOOP_i_13_0_lpi_2_dfm_2 <= STORE_LOOP_i_13_0_lpi_2_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_5_1_2_cse <= 1'b0;
    end
    else if ( core_wen & or_1096_cse & BATCH_LOOP_and_6_tmp & (fsm_output[2]) ) begin
      reg_lfst_exit_STORE_LOOP_lpi_2_dfm_5_1_2_cse <= BATCH_LOOP_acc_1_tmp[4];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm_2_1 <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | or_dcpl_73)) ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm_2_1 <= exit_CONVOLUTION_LOOP_lpi_2_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
          <= 1'b0;
    end
    else if ( core_wen & ((mux_447_nl & BATCH_LOOP_and_6_tmp & (fsm_output[2])) |
        CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1)
        ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
          <= MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_mx0w0,
          CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm,
          CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_for_for_land_2_lpi_2_dfm_st <= 1'b0;
      PADDING_LOOP_for_for_and_psp <= 1'b0;
    end
    else if ( PADDING_LOOP_for_for_aelse_2_and_3_cse ) begin
      PADDING_LOOP_for_for_land_2_lpi_2_dfm_st <= PADDING_LOOP_for_for_land_2_lpi_2_dfm_mx1w0;
      PADDING_LOOP_for_for_and_psp <= PADDING_LOOP_for_for_and_psp_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st <= 1'b0;
      CONVOLUTION_LOOP_for_for_and_psp <= 1'b0;
      reg_CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_ftd_4 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_and_4_cse ) begin
      exit_CONVOLUTION_LOOP_lpi_2_dfm_2_st <= exit_CONVOLUTION_LOOP_lpi_2_dfm_2_mx0w0;
      CONVOLUTION_LOOP_for_for_and_psp <= CONVOLUTION_LOOP_for_for_and_psp_mx1w0;
      reg_CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_ftd_4 <= CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6[0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_PADDING_LOOP_lpi_2_dfm <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | mux_476_nl | (~ BATCH_LOOP_and_6_tmp)))
        ) begin
      exit_PADDING_LOOP_lpi_2_dfm <= exit_PADDING_LOOP_lpi_2_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3 <= 5'b00000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_else_and_836_cse ) begin
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 <= MUX_v_3_2_2((CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0]),
          CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_0, or_tmp_801);
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3 <= MUX_v_5_2_2(CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1,
          CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_7_3, or_tmp_801);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_7_3
          <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_2_0
          <= 3'b000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_if_and_cse ) begin
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_7_3
          <= MUX_v_5_2_2(CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1, CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_7_3,
          or_tmp_805);
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_2_0
          <= MUX_v_3_2_2((CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0]), CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_2_0,
          or_tmp_805);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_1 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_1
          <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1 <= 14'b00000000000000;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_1 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_if_1_and_11_cse ) begin
      CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_1 <= CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1;
      CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_1
          <= CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0];
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1 <= nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1[13:0];
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_1 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_else_mux_973_itm <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_else_mux_972_itm <= 45'b000000000000000000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_else_mux_itm <= 11'b00000000000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_else_and_837_cse ) begin
      CONVOLUTION_LOOP_for_for_for_else_mux_973_itm <= CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_mx0w0;
      CONVOLUTION_LOOP_for_for_for_else_mux_972_itm <= CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_mx0w0;
      CONVOLUTION_LOOP_for_for_for_else_mux_itm <= CONVOLUTION_LOOP_for_for_for_else_mux_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_7_3 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_0 <= 3'b000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_else_and_841_cse ) begin
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_7_3 <= CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_0 <= CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm
          <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | mux_325_cse | (~ BATCH_LOOP_and_6_tmp)))
        ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm
          <= CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st <= 1'b0;
    end
    else if ( core_wen & (~((~ (fsm_output[2])) | or_dcpl_85)) ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_7_3
          <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_2_0
          <= 3'b000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_if_and_833_cse ) begin
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_7_3
          <= CONVOLUTION_LOOP_for_for_for_if_acc_ncse_1;
      CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_2_0
          <= CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1 <= 1'b0;
      lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_1 <= 1'b0;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_2 <= 8'b00000000;
      lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_and_3_cse ) begin
      lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1 <= MUX_s_1_2_2((~ exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4),
          lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2, or_tmp_841);
      lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_1 <= MUX_s_1_2_2((~ exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3),
          lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2, or_tmp_841);
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3 <= MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1,
          exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2, or_tmp_841);
      CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_2 <= MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_3,
          CONVOLUTION_LOOP_for_for_for_y_lpi_2, or_tmp_841);
      lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1 <= MUX_s_1_2_2((~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1),
          lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2, or_tmp_841);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_dfm_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_dfm_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_dfm_1 <= 45'b000000000000000000000000000000000000000000000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_acc_and_1_cse ) begin
      CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_dfm_1 <= MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_0_sva_2,
          CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2, or_tmp_851);
      CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_dfm_1 <= MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_46_sva_2,
          CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2, or_tmp_851);
      CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_dfm_1 <= MUX_v_45_2_2(CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_2,
          CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2, or_tmp_851);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1 <= 8'b00000000;
    end
    else if ( core_wen & (((~ or_tmp_645) & BATCH_LOOP_and_6_tmp & (fsm_output[2]))
        | CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1_mx0c1) ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1 <= MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1,
          CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2, CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_info_index_15_0_lpi_2_dfm <= 16'b0000000000000000;
      PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0 <= 5'b00000;
      CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0 <= 5'b00000;
    end
    else if ( dma_read_info_index_and_itm ) begin
      dma_read_info_index_15_0_lpi_2_dfm <= MUX_v_16_2_2(z_out_6, dma_read_info_index_15_0_lpi_2,
          and_192_nl);
      PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0 <= PADDING_LOOP_chan_5_0_lpi_2_dfm_3_4_0_mx1w0;
      CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0 <= CONVOLUTION_LOOP_fl_5_0_lpi_2_dfm_3_4_0_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_STORE_LOOP_lpi_2_dfm_8_2 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_8_0 <= 1'b0;
      lfst_exit_STORE_LOOP_lpi_2_dfm_8_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2
          <= 1'b0;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_2 <= 1'b0;
      BATCH_LOOP_asn_itm_2 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_else_mux_itm_1 <= 11'b00000000000;
      CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1 <= 45'b000000000000000000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_2 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_2
          <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2 <= 14'b00000000000000;
      CONVOLUTION_LOOP_for_for_for_unequal_tmp_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
          <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
          <= 45'b000000000000000000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1
          <= 1'b0;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2 <= 1'b0;
      STORE_LOOP_equal_tmp_2_2 <= 1'b0;
    end
    else if ( STORE_LOOP_and_726_cse ) begin
      lfst_exit_STORE_LOOP_lpi_2_dfm_8_2 <= STORE_LOOP_STORE_LOOP_or_tmp;
      lfst_exit_STORE_LOOP_lpi_2_dfm_8_0 <= STORE_LOOP_or_2336_tmp;
      lfst_exit_STORE_LOOP_lpi_2_dfm_8_1 <= STORE_LOOP_or_2335_tmp;
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2
          <= CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_2 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_1;
      BATCH_LOOP_asn_itm_2 <= BATCH_LOOP_asn_itm_1;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_2_0 <= CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_1_0;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3 <= MUX_v_5_2_2(CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3,
          CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_7_3,
          and_dcpl_145);
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0 <= MUX_v_3_2_2(CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0,
          CONVOLUTION_LOOP_for_for_for_if_CONVOLUTION_LOOP_for_for_for_if_conc_decb_8_1_sva_1_2_0,
          and_dcpl_145);
      CONVOLUTION_LOOP_for_for_for_else_mux_itm_1 <= MUX_v_11_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_itm_mx0w0,
          CONVOLUTION_LOOP_for_for_for_else_mux_itm, and_dcpl_145);
      CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1 <= MUX_v_45_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_mx0w0,
          CONVOLUTION_LOOP_for_for_for_else_mux_972_itm, and_dcpl_145);
      CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1 <= MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_mx0w0,
          CONVOLUTION_LOOP_for_for_for_else_mux_973_itm, and_dcpl_145);
      CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_2 <= CONVOLUTION_LOOP_for_for_for_if_1_acc_itm_1;
      CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_2
          <= CONVOLUTION_LOOP_for_for_for_if_1_slc_CONVOLUTION_LOOP_for_for_for_if_1_acc_1_sdt_2_0_itm_1;
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2 <= MUX_v_14_2_2(CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1,
          STORE_LOOP_data_asn_itm_1, and_222_nl);
      CONVOLUTION_LOOP_for_for_for_unequal_tmp_1 <= (CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0!=5'b00000);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
          <= CONVOLUTION_LOOP_for_for_for_acc_46_lpi_2_mx1 & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
          <= MUX_v_45_2_2(45'b000000000000000000000000000000000000000000000, CONVOLUTION_LOOP_for_for_for_acc_45_1_lpi_2_mx1,
          CONVOLUTION_LOOP_for_for_for_for_not_2308_nl);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1
          <= CONVOLUTION_LOOP_for_for_for_acc_0_lpi_2_mx1 & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1);
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_2 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_1;
      STORE_LOOP_equal_tmp_2_2 <= STORE_LOOP_equal_tmp_2_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_crt_sva_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      pad_sva <= 8'b00000000;
      dma_read_data_length_sva <= 16'b0000000000000000;
      dma_read_data_length_mul_4_cse_sva <= 16'b0000000000000000;
      n_w_in_acc_psp_sva <= 7'b0000000;
      n_h_in_acc_psp_sva <= 7'b0000000;
      dma_write_data_length_sva <= 16'b0000000000000000;
      n_w_out_lpi_1_dfm <= 8'b00000000;
      n_h_out_lpi_1_dfm <= 8'b00000000;
    end
    else if ( and_986_cse ) begin
      conf_info_crt_sva_231_0 <= conf_info_rsci_idat_mxwt;
      pad_sva <= z_out_5_12_0[7:0];
      dma_read_data_length_sva <= z_out;
      dma_read_data_length_mul_4_cse_sva <= z_out_8_15_0;
      n_w_in_acc_psp_sva <= nl_n_w_in_acc_psp_sva[6:0];
      n_h_in_acc_psp_sva <= nl_n_h_in_acc_psp_sva[6:0];
      dma_write_data_length_sva <= nl_dma_write_data_length_sva[15:0];
      n_w_out_lpi_1_dfm <= MUX_v_8_2_2((z_out_1_8_0[7:0]), asn_3_mx0w1, or_tmp_901);
      n_h_out_lpi_1_dfm <= MUX_v_8_2_2(asn_1_mx0w0, asn_mx0w1, or_tmp_901);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      BATCH_LOOP_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (BATCH_LOOP_stage_v_2_mx0c0 | (BATCH_LOOP_and_4_tmp & (fsm_output[2])))
        ) begin
      BATCH_LOOP_stage_v_2 <= ~ BATCH_LOOP_stage_v_2_mx0c0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      BATCH_LOOP_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (BATCH_LOOP_stage_v_3_mx0c0 | (and_dcpl_128 & (fsm_output[2])))
        ) begin
      BATCH_LOOP_stage_v_3 <= ~ BATCH_LOOP_stage_v_3_mx0c0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_i_lpi_2 <= 16'b0000000000000000;
    end
    else if ( core_wen & ((fsm_output[1]) | LOAD_LOOP_i_lpi_2_mx0c1) ) begin
      LOAD_LOOP_i_lpi_2 <= MUX_v_16_2_2(LOAD_LOOP_i_lpi_2_dfm_2, LOAD_LOOP_i_lpi_2_dfm_2_mx0w0,
          LOAD_LOOP_i_lpi_2_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_for_row_4_0_lpi_2 <= 5'b00000;
      PADDING_LOOP_for_for_col_4_0_lpi_2 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_2 <= 5'b00000;
      STORE_LOOP_i_13_0_lpi_2 <= 14'b00000000000000;
      CONVOLUTION_LOOP_for_for_for_x_lpi_2 <= 8'b00000000;
    end
    else if ( PADDING_LOOP_for_row_and_3_cse ) begin
      PADDING_LOOP_for_row_4_0_lpi_2 <= MUX_v_5_2_2(PADDING_LOOP_for_row_4_0_lpi_2_dfm_5,
          PADDING_LOOP_for_row_4_0_lpi_2_dfm_5_mx0w0, PADDING_LOOP_for_row_and_1_rgt);
      PADDING_LOOP_for_for_col_4_0_lpi_2 <= MUX_v_5_2_2(PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4,
          PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_4_mx0w0, PADDING_LOOP_for_row_and_1_rgt);
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2 <= MUX_v_3_2_2(CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4,
          CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_4_mx0w0, PADDING_LOOP_for_row_and_1_rgt);
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2 <= MUX_v_3_2_2(CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3,
          CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_3_mx0w0, PADDING_LOOP_for_row_and_1_rgt);
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2 <= MUX_v_5_2_2(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5,
          CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_5_mx0w0, PADDING_LOOP_for_row_and_1_rgt);
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_2 <= MUX_v_5_2_2(CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5,
          CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_5_mx0w0, PADDING_LOOP_for_row_and_1_rgt);
      STORE_LOOP_i_13_0_lpi_2 <= MUX_v_14_2_2(STORE_LOOP_i_13_0_lpi_2_dfm_2, STORE_LOOP_i_13_0_lpi_2_dfm_2_mx0w0,
          PADDING_LOOP_for_row_and_1_rgt);
      CONVOLUTION_LOOP_for_for_for_x_lpi_2 <= MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2,
          CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_2_mx0w0, PADDING_LOOP_for_row_and_1_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_PADDING_LOOP_for_lpi_2 <= 1'b0;
      lfst_exit_CONVOLUTION_LOOP_for_lpi_2 <= 1'b0;
    end
    else if ( PADDING_LOOP_for_and_3_cse ) begin
      lfst_exit_PADDING_LOOP_for_lpi_2 <= MUX_s_1_2_2(lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1,
          lfst_exit_PADDING_LOOP_for_lpi_2_dfm_1_mx0w0, fsm_output[2]);
      lfst_exit_CONVOLUTION_LOOP_for_lpi_2 <= MUX_s_1_2_2(lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1,
          lfst_exit_CONVOLUTION_LOOP_for_lpi_2_dfm_1_mx0w0, fsm_output[2]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2 <= 1'b0;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2 <= 1'b0;
      lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2 <= 1'b0;
      lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_for_and_12_cse ) begin
      lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2 <= MUX_s_1_2_2(lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1,
          (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1), fsm_output[2]);
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2 <= MUX_s_1_2_2(exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3,
          exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_mx0w1, fsm_output[2]);
      lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2 <= MUX_s_1_2_2(lfst_exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_1,
          (~ exit_CONVOLUTION_LOOP_for_for_for_lpi_2_dfm_3), fsm_output[2]);
      lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2 <= MUX_s_1_2_2(lfst_exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_1,
          (~ exit_CONVOLUTION_LOOP_for_for_lpi_2_dfm_4), fsm_output[2]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      BATCH_LOOP_stage_0_3 <= 1'b0;
    end
    else if ( core_wen & ((fsm_output[1]) | ((and_dcpl_128 | BATCH_LOOP_and_4_tmp)
        & (fsm_output[2]))) ) begin
      BATCH_LOOP_stage_0_3 <= BATCH_LOOP_stage_0_2 & (~ (fsm_output[1]));
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_y_lpi_2 <= 8'b00000000;
    end
    else if ( core_wen & ((~ (fsm_output[2])) | CONVOLUTION_LOOP_for_for_for_y_and_4_rgt)
        ) begin
      CONVOLUTION_LOOP_for_for_for_y_lpi_2 <= MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_2,
          CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_3, CONVOLUTION_LOOP_for_for_for_y_and_4_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2 <= 8'b00000000;
    end
    else if ( core_wen & ((~ (fsm_output[2])) | CONVOLUTION_LOOP_for_for_for_y_and_2_rgt)
        ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2 <= MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_2_dfm_1,
          CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1, CONVOLUTION_LOOP_for_for_for_y_and_2_rgt);
    end
  end
  assign mux_525_nl = MUX_s_1_2_2(or_tmp_372, and_830_cse, STORE_LOOP_or_2336_tmp);
  assign mux_526_nl = MUX_s_1_2_2(mux_525_nl, exitL_exit_STORE_LOOP_sva, or_214_cse);
  assign mux_528_nl = MUX_s_1_2_2((~ BATCH_LOOP_stage_v), mux_tmp_355, BATCH_LOOP_and_6_tmp);
  assign nor_246_nl = ~(or_tmp_369 | (~(lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2 & or_tmp_16)));
  assign mux_534_nl = MUX_s_1_2_2(or_tmp_16, nor_246_nl, and_dcpl_32);
  assign or_779_nl = or_tmp_284 | and_830_cse | nand_tmp_57;
  assign or_776_nl = or_81_cse | nand_tmp_57;
  assign mux_537_nl = MUX_s_1_2_2(or_779_nl, or_776_nl, or_214_cse);
  assign or_780_nl = mux_537_nl | (BATCH_LOOP_acc_1_tmp[4]) | (~ BATCH_LOOP_and_6_tmp);
  assign STORE_LOOP_mux_37_nl = MUX_v_4_2_2((BATCH_LOOP_acc_1_tmp[3:0]), BATCH_LOOP_b_4_0_sva_3_0,
      or_780_nl);
  assign PADDING_LOOP_for_for_aelse_mux_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_1, BATCH_LOOP_stage_0,
      BATCH_LOOP_and_6_tmp);
  assign nor_379_nl = ~(BATCH_LOOP_and_4_tmp | BATCH_LOOP_and_6_tmp);
  assign BATCH_LOOP_mux_5_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_1, BATCH_LOOP_stage_0_2,
      nor_379_nl);
  assign or_6_nl = plm_f_data_rsci_bawt | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2;
  assign mux_531_nl = MUX_s_1_2_2(not_tmp_312, or_2_cse, or_6_nl);
  assign or_1_nl = plm_in_data_rsci_bawt | lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_2;
  assign mux_530_nl = MUX_s_1_2_2(not_tmp_312, or_2_cse, or_1_nl);
  assign mux_532_nl = MUX_s_1_2_2(mux_531_nl, mux_530_nl, lfst_exit_STORE_LOOP_lpi_2_dfm_st_2_0);
  assign nand_65_nl = ~(BATCH_LOOP_stage_0_3 & BATCH_LOOP_stage_v_2 & mux_532_nl);
  assign nand_66_nl = ~((lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_0 | lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_1
      | (~ lfst_exit_STORE_LOOP_lpi_2_dfm_st_3_2) | (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_3_st_3)
      | (~ CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3)
      | plm_out_data_rsci_bawt) & BATCH_LOOP_stage_0_4 & or_2_cse);
  assign mux_533_nl = MUX_s_1_2_2(nand_65_nl, nand_66_nl, BATCH_LOOP_stage_v_3);
  assign BATCH_LOOP_mux_6_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_3, BATCH_LOOP_stage_0_4,
      mux_533_nl);
  assign mux_331_nl = MUX_s_1_2_2(nand_tmp_29, or_tmp_314, or_214_cse);
  assign PADDING_LOOP_for_for_index_in_mul_2_nl = conv_u2u_13_13(PADDING_LOOP_for_row_4_0_lpi_2
      * ({n_h_in_acc_psp_sva , (conf_info_crt_sva_231_0[160])}));
  assign nl_PADDING_LOOP_for_for_index_in_acc_2_nl = PADDING_LOOP_for_for_index_in_mul_2_nl
      + conv_u2u_5_13(PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5);
  assign PADDING_LOOP_for_for_index_in_acc_2_nl = nl_PADDING_LOOP_for_for_index_in_acc_2_nl[12:0];
  assign PADDING_LOOP_for_for_index_in_mul_1_nl = conv_u2u_13_13(PADDING_LOOP_chan_5_0_lpi_2_4_0
      * ({n_w_in_acc_psp_sva , (conf_info_crt_sva_231_0[192])}));
  assign nl_PADDING_LOOP_for_for_index_in_mul_nl = PADDING_LOOP_for_for_index_in_mul_1_nl
      * ({n_h_in_acc_psp_sva , (conf_info_crt_sva_231_0[160])});
  assign PADDING_LOOP_for_for_index_in_mul_nl = nl_PADDING_LOOP_for_for_index_in_mul_nl[13:0];
  assign nl_PADDING_LOOP_for_for_index_in_acc_itm_1  = conv_u2u_13_14(PADDING_LOOP_for_for_index_in_acc_2_nl)
      + PADDING_LOOP_for_for_index_in_mul_nl;
  assign and_764_nl = nor_tmp_142 & (~ or_tmp_444);
  assign nor_232_nl = ~(or_131_cse | (~ or_tmp_440));
  assign mux_378_nl = MUX_s_1_2_2(and_764_nl, nor_232_nl, or_214_cse);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl = CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_mx0
      * ({n_w_in_acc_psp_sva , (conf_info_crt_sva_231_0[192])});
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl
      + conv_u2u_8_14(CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_mx0);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl = ({n_w_in_acc_psp_sva
      , (conf_info_crt_sva_231_0[192])}) * ({n_h_in_acc_psp_sva , (conf_info_crt_sva_231_0[160])});
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl
      * CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1;
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1  = CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl
      + CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl;
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl = z_out_5_12_0 * (conf_info_crt_sva_231_0[103:96]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl[15:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_5_nl = conv_u2u_11_11(CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_2_dfm_4
      * (conf_info_crt_sva_231_0[103:96]));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_5_nl
      + conv_u2u_3_11(CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_2_dfm_5);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl[10:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl
      + conv_u2u_11_16(CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl[15:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1  = CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl
      + z_out_9_15_0;
  assign and_762_nl = (~((~ BATCH_LOOP_and_4_tmp) | BATCH_LOOP_asn_itm_1 | STORE_LOOP_or_2335_tmp
      | STORE_LOOP_or_2336_tmp | (~ STORE_LOOP_STORE_LOOP_or_tmp))) & not_tmp_258;
  assign or_603_nl = (~ CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp) | (operator_8_false_4_acc_tmp[8:3]!=6'b000000)
      | (~ or_tmp_509);
  assign mux_444_nl = MUX_s_1_2_2((~ or_tmp_509), or_603_nl, operator_8_false_8_acc_itm_3_1);
  assign nand_49_nl = ~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & (~(nor_229_cse
      | (operator_8_false_4_acc_tmp[8:3]!=6'b000000) | (~ or_tmp_509))));
  assign mux_445_nl = MUX_s_1_2_2(mux_444_nl, nand_49_nl, operator_8_false_9_acc_itm_3_1);
  assign nor_227_nl = ~(exitL_exit_STORE_LOOP_sva | mux_445_nl);
  assign and_763_nl = (~(STORE_LOOP_or_2335_tmp | STORE_LOOP_or_2336_tmp | (~ STORE_LOOP_STORE_LOOP_or_tmp)))
      & not_tmp_258;
  assign nor_230_nl = ~(exitL_exit_STORE_LOOP_sva | mux_tmp_435);
  assign mux_443_nl = MUX_s_1_2_2(and_763_nl, nor_230_nl, BATCH_LOOP_asn_itm_1);
  assign mux_446_nl = MUX_s_1_2_2(nor_227_nl, mux_443_nl, BATCH_LOOP_and_4_tmp);
  assign nor_187_nl = ~(lfst_exit_STORE_LOOP_lpi_2_1 | lfst_exit_STORE_LOOP_lpi_2_0
      | (~ lfst_exit_STORE_LOOP_lpi_2_2));
  assign mux_447_nl = MUX_s_1_2_2(and_762_nl, mux_446_nl, nor_187_nl);
  assign or_636_nl = (~ PADDING_LOOP_for_if_equal_tmp) | (operator_8_false_2_acc_tmp[8:5]!=4'b0000)
      | mux_tmp_357;
  assign mux_476_nl = MUX_s_1_2_2(mux_tmp_357, or_636_nl, operator_8_false_2_acc_itm_4_1);
  assign CONVOLUTION_LOOP_for_for_for_index_out_mul_2_nl = conv_u2u_13_13(CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6
      * n_w_out_lpi_1_dfm);
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl = CONVOLUTION_LOOP_for_for_for_index_out_mul_2_nl
      + conv_u2u_5_13(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_2_dfm_6);
  assign CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl = nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl[12:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl = n_w_out_lpi_1_dfm *
      n_h_out_lpi_1_dfm;
  assign CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl = nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_nl = CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl
      * CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0;
  assign CONVOLUTION_LOOP_for_for_for_index_out_mul_nl = nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1  = conv_u2u_13_14(CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl)
      + CONVOLUTION_LOOP_for_for_for_index_out_mul_nl;
  assign and_192_nl = (~ mux_tmp_354) & BATCH_LOOP_and_6_tmp;
  assign and_222_nl = BATCH_LOOP_and_4_tmp & reg_lfst_exit_STORE_LOOP_lpi_2_dfm_1_0_cse;
  assign CONVOLUTION_LOOP_for_for_for_for_not_2308_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_2_dfm_1;
  assign nl_n_w_in_acc_psp_sva  = (conf_info_rsci_idat_mxwt[199:193]) + (z_out_5_12_0[6:0]);
  assign nl_n_h_in_acc_psp_sva  = (conf_info_rsci_idat_mxwt[167:161]) + (z_out_5_12_0[6:0]);
  assign nl_dma_write_data_length_sva  = z_out_9_15_0 * (conf_info_rsci_idat_mxwt[71:64]);
  assign BATCH_LOOP_mux_10_nl = MUX_v_16_2_2(z_out_8_15_0, z_out_6, fsm_output[1]);
  assign nl_BATCH_LOOP_mul_3_nl = dma_write_data_length_sva * BATCH_LOOP_b_4_0_sva_3_0;
  assign BATCH_LOOP_mul_3_nl = nl_BATCH_LOOP_mul_3_nl[15:0];
  assign nl_dma_read_data_length_mul_5_nl = (z_out_7[15:0]) * (conf_info_rsci_idat_mxwt[71:64]);
  assign dma_read_data_length_mul_5_nl = nl_dma_read_data_length_mul_5_nl[15:0];
  assign BATCH_LOOP_mux_11_nl = MUX_v_16_2_2(BATCH_LOOP_mul_3_nl, dma_read_data_length_mul_5_nl,
      fsm_output[1]);
  assign nl_z_out = BATCH_LOOP_mux_10_nl + BATCH_LOOP_mux_11_nl;
  assign z_out = nl_z_out[15:0];
  assign operator_42_true_mux_2_nl = MUX_v_9_2_2((signext_9_8(else_acc_psp_sva_1[8:1])),
      ({4'b1000 , PADDING_LOOP_for_for_col_4_0_lpi_2_dfm_5}), fsm_output[2]);
  assign operator_42_true_and_1_nl = (else_acc_psp_sva_1[10]) & (else_acc_psp_sva_1[0]);
  assign operator_42_true_mux_3_nl = MUX_v_8_2_2(({7'b0000000 , operator_42_true_and_1_nl}),
      (~ pad_sva), fsm_output[2]);
  assign nl_acc_1_nl = ({operator_42_true_mux_2_nl , 1'b1}) + conv_u2u_9_10({operator_42_true_mux_3_nl
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[9:0];
  assign z_out_1_8_0 = readslicef_10_9_1(acc_1_nl);
  assign nl_PADDING_LOOP_for_for_aelse_2_acc_2_nl = conv_u2u_8_9({(~ n_w_in_acc_psp_sva)
      , (~ (conf_info_crt_sva_231_0[192]))}) + conv_u2u_8_9(pad_sva) + 9'b000000001;
  assign PADDING_LOOP_for_for_aelse_2_acc_2_nl = nl_PADDING_LOOP_for_for_aelse_2_acc_2_nl[8:0];
  assign else_mux_2_nl = MUX_v_9_2_2(({(z_out_5_12_0[7:0]) , 1'b0}), PADDING_LOOP_for_for_aelse_2_acc_2_nl,
      fsm_output[2]);
  assign else_or_1_nl = (fsm_output[2:1]!=2'b10);
  assign else_else_nor_1_nl = ~(MUX_v_3_2_2((conf_info_rsci_idat_mxwt[103:101]),
      3'b111, (fsm_output[2])));
  assign else_mux_3_nl = MUX_v_5_2_2((~ (conf_info_rsci_idat_mxwt[100:96])), PADDING_LOOP_for_row_4_0_lpi_2,
      fsm_output[2]);
  assign nl_acc_2_nl = conv_u2u_10_11({else_mux_2_nl , else_or_1_nl}) + conv_s2u_10_11({(fsm_output[2])
      , else_else_nor_1_nl , else_mux_3_nl , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[10:0];
  assign z_out_2 = readslicef_11_10_1(acc_2_nl);
  assign pad_pad_pad_nor_1_nl = ~(MUX_v_3_2_2((conf_info_rsci_idat_mxwt[199:197]),
      3'b111, (fsm_output[2])));
  assign pad_mux_5_nl = MUX_v_5_2_2((~ (conf_info_rsci_idat_mxwt[196:192])), PADDING_LOOP_for_row_4_0_lpi_2,
      fsm_output[2]);
  assign pad_mux_6_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[103:96]), (~ pad_sva),
      fsm_output[2]);
  assign nl_acc_3_nl = ({1'b1 , pad_pad_pad_nor_1_nl , pad_mux_5_nl , 1'b1}) + conv_u2u_9_10({pad_mux_6_nl
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[9:0];
  assign z_out_3 = readslicef_10_9_1(acc_3_nl);
  assign operator_8_false_mux_1_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[199:192]),
      (conf_info_crt_sva_231_0[135:128]), fsm_output[2]);
  assign nl_z_out_4 = conv_u2u_8_9(operator_8_false_mux_1_nl) + 9'b111111111;
  assign z_out_4 = nl_z_out_4[8:0];
  assign operator_43_true_and_1_nl = (z_out_12[16]) & (z_out_12[0]);
  assign nl_operator_43_true_operator_43_true_acc_1_nl = (z_out_12[8:1]) + conv_u2s_1_8(operator_43_true_and_1_nl);
  assign operator_43_true_operator_43_true_acc_1_nl = nl_operator_43_true_operator_43_true_acc_1_nl[7:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_10_nl = MUX_v_8_2_2(({3'b000 ,
      CONVOLUTION_LOOP_for_k_5_0_lpi_2_4_0_mx1}), operator_43_true_operator_43_true_acc_1_nl,
      fsm_output[1]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_11_nl = MUX_v_8_2_2((conf_info_crt_sva_231_0[103:96]),
      (conf_info_rsci_idat_mxwt[39:32]), fsm_output[1]);
  assign nl_z_out_5_12_0 = CONVOLUTION_LOOP_for_for_for_for_for_mux_10_nl * CONVOLUTION_LOOP_for_for_for_for_for_mux_11_nl;
  assign z_out_5_12_0 = nl_z_out_5_12_0[12:0];
  assign dma_read_data_length_mux_8_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[135:128]),
      ({4'b0000 , BATCH_LOOP_b_4_0_sva_3_0}), fsm_output[2]);
  assign dma_read_data_length_mux_9_nl = MUX_v_16_2_2((z_out_10[15:0]), dma_read_data_length_sva,
      fsm_output[2]);
  assign nl_z_out_6 = dma_read_data_length_mux_8_nl * dma_read_data_length_mux_9_nl;
  assign z_out_6 = nl_z_out_6[15:0];
  assign dma_read_data_length_mux_10_nl = MUX_v_32_2_2(({16'b0000000000000000 , z_out_8_15_0}),
      plm_f_data_rsci_q_d_mxwt, fsm_output[2]);
  assign dma_read_data_length_mux_11_nl = MUX_v_32_2_2(({24'b000000000000000000000000
      , (conf_info_rsci_idat_mxwt[135:128])}), plm_in_data_rsci_q_d_mxwt, fsm_output[2]);
  assign z_out_7 = conv_u2u_64_64($signed(dma_read_data_length_mux_10_nl) * $signed(dma_read_data_length_mux_11_nl));
  assign BATCH_LOOP_mux_12_nl = MUX_v_8_2_2((conf_info_crt_sva_231_0[231:224]), (conf_info_rsci_idat_mxwt[103:96]),
      fsm_output[1]);
  assign BATCH_LOOP_mux_13_nl = MUX_v_16_2_2(dma_read_data_length_sva, ({8'b00000000
      , (conf_info_rsci_idat_mxwt[103:96])}), fsm_output[1]);
  assign nl_z_out_8_15_0 = $signed(conv_u2s_8_9(BATCH_LOOP_mux_12_nl)) * $signed(BATCH_LOOP_mux_13_nl);
  assign z_out_8_15_0 = nl_z_out_8_15_0[15:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_14_nl = (~ and_dcpl_138) & (fsm_output[1]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_mux1h_2_nl
      = MUX1HOT_v_8_3_2((conf_info_crt_sva_231_0[135:128]), asn_1_mx0w0, asn_mx0w1,
      {(~ (fsm_output[1])) , CONVOLUTION_LOOP_for_for_for_for_for_and_14_nl , or_tmp_901});
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_11_nl = conv_u2u_13_13(CONVOLUTION_LOOP_fl_5_0_lpi_2_4_0
      * (conf_info_crt_sva_231_0[103:96]));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_10_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_11_nl
      * (conf_info_crt_sva_231_0[103:96]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_10_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_10_nl[15:0];
  assign mux_562_nl = MUX_v_8_2_2((z_out_1_8_0[7:0]), asn_3_mx0w1, and_dcpl_138);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_12_nl = MUX_v_16_2_2(CONVOLUTION_LOOP_for_for_for_for_for_mul_10_nl,
      ({8'b00000000 , mux_562_nl}), fsm_output[1]);
  assign nl_z_out_9_15_0 = $signed(conv_u2s_8_9(CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_mux1h_2_nl))
      * $signed(CONVOLUTION_LOOP_for_for_for_for_for_mux_12_nl);
  assign z_out_9_15_0 = nl_z_out_9_15_0[15:0];
  assign dma_read_data_length_mux_12_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[167:160]),
      (conf_info_crt_sva_231_0[71:64]), fsm_output[2]);
  assign LOAD_LOOP_mul_2_nl = conv_u2u_24_24(dma_read_data_length_mul_4_cse_sva *
      (conf_info_crt_sva_231_0[135:128]));
  assign dma_read_data_length_mux_13_nl = MUX_v_24_2_2(({16'b0000000000000000 , (conf_info_rsci_idat_mxwt[199:192])}),
      LOAD_LOOP_mul_2_nl, fsm_output[2]);
  assign z_out_10 = conv_u2u_32_32(dma_read_data_length_mux_12_nl * dma_read_data_length_mux_13_nl);
  assign pad_mux_7_nl = MUX_v_8_2_2((conf_info_rsci_idat_mxwt[7:0]), ({3'b000 , CONVOLUTION_LOOP_for_for_i_4_0_lpi_2_dfm_6}),
      fsm_output[2]);
  assign pad_mux_8_nl = MUX_v_9_2_2(z_out_4, ({1'b0 , (conf_info_crt_sva_231_0[7:0])}),
      fsm_output[2]);
  assign nl_z_out_11_16_0 = $signed(conv_u2s_8_9(pad_mux_7_nl)) * $signed(pad_mux_8_nl);
  assign z_out_11_16_0 = nl_z_out_11_16_0[16:0];
  assign LOAD_LOOP_mux_2_nl = MUX_v_17_2_2(({1'b0 , LOAD_LOOP_i_lpi_2_mx1}), z_out_11_16_0,
      fsm_output[1]);
  assign LOAD_LOOP_mux_3_nl = MUX_v_9_2_2(9'b000000001, z_out_3, fsm_output[1]);
  assign nl_z_out_12 = LOAD_LOOP_mux_2_nl + conv_s2u_9_17(LOAD_LOOP_mux_3_nl);
  assign z_out_12 = nl_z_out_12[16:0];
  assign and_987_nl = or_1062_cse & operator_8_false_9_acc_itm_3_1 & (fsm_output[2]);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2951_nl = MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_x_lpi_2_dfm_mx0,
      CONVOLUTION_LOOP_for_for_for_y_lpi_2_dfm_mx0, and_987_nl);
  assign nl_z_out_13 = CONVOLUTION_LOOP_for_for_for_for_mux_2951_nl + 8'b00000001;
  assign z_out_13 = nl_z_out_13[7:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [13:0] MUX1HOT_v_14_3_2;
    input [13:0] input_2;
    input [13:0] input_1;
    input [13:0] input_0;
    input [2:0] sel;
    reg [13:0] result;
  begin
    result = input_0 & {14{sel[0]}};
    result = result | ( input_1 & {14{sel[1]}});
    result = result | ( input_2 & {14{sel[2]}});
    MUX1HOT_v_14_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [44:0] MUX1HOT_v_45_3_2;
    input [44:0] input_2;
    input [44:0] input_1;
    input [44:0] input_0;
    input [2:0] sel;
    reg [44:0] result;
  begin
    result = input_0 & {45{sel[0]}};
    result = result | ( input_1 & {45{sel[1]}});
    result = result | ( input_2 & {45{sel[2]}});
    MUX1HOT_v_45_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_324_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] input_2;
    input [0:0] input_3;
    input [0:0] input_4;
    input [0:0] input_5;
    input [0:0] input_6;
    input [0:0] input_7;
    input [0:0] input_8;
    input [0:0] input_9;
    input [0:0] input_10;
    input [0:0] input_11;
    input [0:0] input_12;
    input [0:0] input_13;
    input [0:0] input_14;
    input [0:0] input_15;
    input [0:0] input_16;
    input [0:0] input_17;
    input [0:0] input_18;
    input [0:0] input_19;
    input [0:0] input_20;
    input [0:0] input_21;
    input [0:0] input_22;
    input [0:0] input_23;
    input [0:0] input_24;
    input [0:0] input_25;
    input [0:0] input_26;
    input [0:0] input_27;
    input [0:0] input_28;
    input [0:0] input_29;
    input [0:0] input_30;
    input [0:0] input_31;
    input [0:0] input_32;
    input [0:0] input_33;
    input [0:0] input_34;
    input [0:0] input_35;
    input [0:0] input_36;
    input [0:0] input_37;
    input [0:0] input_38;
    input [0:0] input_39;
    input [0:0] input_40;
    input [0:0] input_41;
    input [0:0] input_42;
    input [0:0] input_43;
    input [0:0] input_44;
    input [0:0] input_45;
    input [0:0] input_46;
    input [0:0] input_47;
    input [0:0] input_48;
    input [0:0] input_49;
    input [0:0] input_50;
    input [0:0] input_51;
    input [0:0] input_52;
    input [0:0] input_53;
    input [0:0] input_54;
    input [0:0] input_55;
    input [0:0] input_56;
    input [0:0] input_57;
    input [0:0] input_58;
    input [0:0] input_59;
    input [0:0] input_60;
    input [0:0] input_61;
    input [0:0] input_62;
    input [0:0] input_63;
    input [0:0] input_64;
    input [0:0] input_65;
    input [0:0] input_66;
    input [0:0] input_67;
    input [0:0] input_68;
    input [0:0] input_69;
    input [0:0] input_70;
    input [0:0] input_71;
    input [0:0] input_72;
    input [0:0] input_73;
    input [0:0] input_74;
    input [0:0] input_75;
    input [0:0] input_76;
    input [0:0] input_77;
    input [0:0] input_78;
    input [0:0] input_79;
    input [0:0] input_80;
    input [0:0] input_81;
    input [0:0] input_82;
    input [0:0] input_83;
    input [0:0] input_84;
    input [0:0] input_85;
    input [0:0] input_86;
    input [0:0] input_87;
    input [0:0] input_88;
    input [0:0] input_89;
    input [0:0] input_90;
    input [0:0] input_91;
    input [0:0] input_92;
    input [0:0] input_93;
    input [0:0] input_94;
    input [0:0] input_95;
    input [0:0] input_96;
    input [0:0] input_97;
    input [0:0] input_98;
    input [0:0] input_99;
    input [0:0] input_100;
    input [0:0] input_101;
    input [0:0] input_102;
    input [0:0] input_103;
    input [0:0] input_104;
    input [0:0] input_105;
    input [0:0] input_106;
    input [0:0] input_107;
    input [0:0] input_108;
    input [0:0] input_109;
    input [0:0] input_110;
    input [0:0] input_111;
    input [0:0] input_112;
    input [0:0] input_113;
    input [0:0] input_114;
    input [0:0] input_115;
    input [0:0] input_116;
    input [0:0] input_117;
    input [0:0] input_118;
    input [0:0] input_119;
    input [0:0] input_120;
    input [0:0] input_121;
    input [0:0] input_122;
    input [0:0] input_123;
    input [0:0] input_124;
    input [0:0] input_125;
    input [0:0] input_126;
    input [0:0] input_127;
    input [0:0] input_128;
    input [0:0] input_129;
    input [0:0] input_130;
    input [0:0] input_131;
    input [0:0] input_132;
    input [0:0] input_133;
    input [0:0] input_134;
    input [0:0] input_135;
    input [0:0] input_136;
    input [0:0] input_137;
    input [0:0] input_138;
    input [0:0] input_139;
    input [0:0] input_140;
    input [0:0] input_141;
    input [0:0] input_142;
    input [0:0] input_143;
    input [0:0] input_144;
    input [0:0] input_145;
    input [0:0] input_146;
    input [0:0] input_147;
    input [0:0] input_148;
    input [0:0] input_149;
    input [0:0] input_150;
    input [0:0] input_151;
    input [0:0] input_152;
    input [0:0] input_153;
    input [0:0] input_154;
    input [0:0] input_155;
    input [0:0] input_156;
    input [0:0] input_157;
    input [0:0] input_158;
    input [0:0] input_159;
    input [0:0] input_160;
    input [0:0] input_161;
    input [0:0] input_162;
    input [0:0] input_163;
    input [0:0] input_164;
    input [0:0] input_165;
    input [0:0] input_166;
    input [0:0] input_167;
    input [0:0] input_168;
    input [0:0] input_169;
    input [0:0] input_170;
    input [0:0] input_171;
    input [0:0] input_172;
    input [0:0] input_173;
    input [0:0] input_174;
    input [0:0] input_175;
    input [0:0] input_176;
    input [0:0] input_177;
    input [0:0] input_178;
    input [0:0] input_179;
    input [0:0] input_180;
    input [0:0] input_181;
    input [0:0] input_182;
    input [0:0] input_183;
    input [0:0] input_184;
    input [0:0] input_185;
    input [0:0] input_186;
    input [0:0] input_187;
    input [0:0] input_188;
    input [0:0] input_189;
    input [0:0] input_190;
    input [0:0] input_191;
    input [0:0] input_192;
    input [0:0] input_193;
    input [0:0] input_194;
    input [0:0] input_195;
    input [0:0] input_196;
    input [0:0] input_197;
    input [0:0] input_198;
    input [0:0] input_199;
    input [0:0] input_200;
    input [0:0] input_201;
    input [0:0] input_202;
    input [0:0] input_203;
    input [0:0] input_204;
    input [0:0] input_205;
    input [0:0] input_206;
    input [0:0] input_207;
    input [0:0] input_208;
    input [0:0] input_209;
    input [0:0] input_210;
    input [0:0] input_211;
    input [0:0] input_212;
    input [0:0] input_213;
    input [0:0] input_214;
    input [0:0] input_215;
    input [0:0] input_216;
    input [0:0] input_217;
    input [0:0] input_218;
    input [0:0] input_219;
    input [0:0] input_220;
    input [0:0] input_221;
    input [0:0] input_222;
    input [0:0] input_223;
    input [0:0] input_224;
    input [0:0] input_225;
    input [0:0] input_226;
    input [0:0] input_227;
    input [0:0] input_228;
    input [0:0] input_229;
    input [0:0] input_230;
    input [0:0] input_231;
    input [0:0] input_232;
    input [0:0] input_233;
    input [0:0] input_234;
    input [0:0] input_235;
    input [0:0] input_236;
    input [0:0] input_237;
    input [0:0] input_238;
    input [0:0] input_239;
    input [0:0] input_240;
    input [0:0] input_241;
    input [0:0] input_242;
    input [0:0] input_243;
    input [0:0] input_244;
    input [0:0] input_245;
    input [0:0] input_246;
    input [0:0] input_247;
    input [0:0] input_248;
    input [0:0] input_249;
    input [0:0] input_250;
    input [0:0] input_251;
    input [0:0] input_252;
    input [0:0] input_253;
    input [0:0] input_254;
    input [0:0] input_255;
    input [0:0] input_256;
    input [0:0] input_257;
    input [0:0] input_258;
    input [0:0] input_259;
    input [0:0] input_260;
    input [0:0] input_261;
    input [0:0] input_262;
    input [0:0] input_263;
    input [0:0] input_264;
    input [0:0] input_265;
    input [0:0] input_266;
    input [0:0] input_267;
    input [0:0] input_268;
    input [0:0] input_269;
    input [0:0] input_270;
    input [0:0] input_271;
    input [0:0] input_272;
    input [0:0] input_273;
    input [0:0] input_274;
    input [0:0] input_275;
    input [0:0] input_276;
    input [0:0] input_277;
    input [0:0] input_278;
    input [0:0] input_279;
    input [0:0] input_280;
    input [0:0] input_281;
    input [0:0] input_282;
    input [0:0] input_283;
    input [0:0] input_284;
    input [0:0] input_285;
    input [0:0] input_286;
    input [0:0] input_287;
    input [0:0] input_288;
    input [0:0] input_289;
    input [0:0] input_290;
    input [0:0] input_291;
    input [0:0] input_292;
    input [0:0] input_293;
    input [0:0] input_294;
    input [0:0] input_295;
    input [0:0] input_296;
    input [0:0] input_297;
    input [0:0] input_298;
    input [0:0] input_299;
    input [0:0] input_300;
    input [0:0] input_301;
    input [0:0] input_302;
    input [0:0] input_303;
    input [0:0] input_304;
    input [0:0] input_305;
    input [0:0] input_306;
    input [0:0] input_307;
    input [0:0] input_308;
    input [0:0] input_309;
    input [0:0] input_310;
    input [0:0] input_311;
    input [0:0] input_312;
    input [0:0] input_313;
    input [0:0] input_314;
    input [0:0] input_315;
    input [0:0] input_316;
    input [0:0] input_317;
    input [0:0] input_318;
    input [0:0] input_319;
    input [0:0] input_320;
    input [0:0] input_321;
    input [0:0] input_322;
    input [0:0] input_323;
    input [8:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_s_1_324_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_324_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [10:0] input_8;
    input [10:0] input_9;
    input [10:0] input_10;
    input [10:0] input_11;
    input [10:0] input_12;
    input [10:0] input_13;
    input [10:0] input_14;
    input [10:0] input_15;
    input [10:0] input_16;
    input [10:0] input_17;
    input [10:0] input_18;
    input [10:0] input_19;
    input [10:0] input_20;
    input [10:0] input_21;
    input [10:0] input_22;
    input [10:0] input_23;
    input [10:0] input_24;
    input [10:0] input_25;
    input [10:0] input_26;
    input [10:0] input_27;
    input [10:0] input_28;
    input [10:0] input_29;
    input [10:0] input_30;
    input [10:0] input_31;
    input [10:0] input_32;
    input [10:0] input_33;
    input [10:0] input_34;
    input [10:0] input_35;
    input [10:0] input_36;
    input [10:0] input_37;
    input [10:0] input_38;
    input [10:0] input_39;
    input [10:0] input_40;
    input [10:0] input_41;
    input [10:0] input_42;
    input [10:0] input_43;
    input [10:0] input_44;
    input [10:0] input_45;
    input [10:0] input_46;
    input [10:0] input_47;
    input [10:0] input_48;
    input [10:0] input_49;
    input [10:0] input_50;
    input [10:0] input_51;
    input [10:0] input_52;
    input [10:0] input_53;
    input [10:0] input_54;
    input [10:0] input_55;
    input [10:0] input_56;
    input [10:0] input_57;
    input [10:0] input_58;
    input [10:0] input_59;
    input [10:0] input_60;
    input [10:0] input_61;
    input [10:0] input_62;
    input [10:0] input_63;
    input [10:0] input_64;
    input [10:0] input_65;
    input [10:0] input_66;
    input [10:0] input_67;
    input [10:0] input_68;
    input [10:0] input_69;
    input [10:0] input_70;
    input [10:0] input_71;
    input [10:0] input_72;
    input [10:0] input_73;
    input [10:0] input_74;
    input [10:0] input_75;
    input [10:0] input_76;
    input [10:0] input_77;
    input [10:0] input_78;
    input [10:0] input_79;
    input [10:0] input_80;
    input [10:0] input_81;
    input [10:0] input_82;
    input [10:0] input_83;
    input [10:0] input_84;
    input [10:0] input_85;
    input [10:0] input_86;
    input [10:0] input_87;
    input [10:0] input_88;
    input [10:0] input_89;
    input [10:0] input_90;
    input [10:0] input_91;
    input [10:0] input_92;
    input [10:0] input_93;
    input [10:0] input_94;
    input [10:0] input_95;
    input [10:0] input_96;
    input [10:0] input_97;
    input [10:0] input_98;
    input [10:0] input_99;
    input [10:0] input_100;
    input [10:0] input_101;
    input [10:0] input_102;
    input [10:0] input_103;
    input [10:0] input_104;
    input [10:0] input_105;
    input [10:0] input_106;
    input [10:0] input_107;
    input [10:0] input_108;
    input [10:0] input_109;
    input [10:0] input_110;
    input [10:0] input_111;
    input [10:0] input_112;
    input [10:0] input_113;
    input [10:0] input_114;
    input [10:0] input_115;
    input [10:0] input_116;
    input [10:0] input_117;
    input [10:0] input_118;
    input [10:0] input_119;
    input [10:0] input_120;
    input [10:0] input_121;
    input [10:0] input_122;
    input [10:0] input_123;
    input [10:0] input_124;
    input [10:0] input_125;
    input [10:0] input_126;
    input [10:0] input_127;
    input [10:0] input_128;
    input [10:0] input_129;
    input [10:0] input_130;
    input [10:0] input_131;
    input [10:0] input_132;
    input [10:0] input_133;
    input [10:0] input_134;
    input [10:0] input_135;
    input [10:0] input_136;
    input [10:0] input_137;
    input [10:0] input_138;
    input [10:0] input_139;
    input [10:0] input_140;
    input [10:0] input_141;
    input [10:0] input_142;
    input [10:0] input_143;
    input [10:0] input_144;
    input [10:0] input_145;
    input [10:0] input_146;
    input [10:0] input_147;
    input [10:0] input_148;
    input [10:0] input_149;
    input [10:0] input_150;
    input [10:0] input_151;
    input [10:0] input_152;
    input [10:0] input_153;
    input [10:0] input_154;
    input [10:0] input_155;
    input [10:0] input_156;
    input [10:0] input_157;
    input [10:0] input_158;
    input [10:0] input_159;
    input [10:0] input_160;
    input [10:0] input_161;
    input [10:0] input_162;
    input [10:0] input_163;
    input [10:0] input_164;
    input [10:0] input_165;
    input [10:0] input_166;
    input [10:0] input_167;
    input [10:0] input_168;
    input [10:0] input_169;
    input [10:0] input_170;
    input [10:0] input_171;
    input [10:0] input_172;
    input [10:0] input_173;
    input [10:0] input_174;
    input [10:0] input_175;
    input [10:0] input_176;
    input [10:0] input_177;
    input [10:0] input_178;
    input [10:0] input_179;
    input [10:0] input_180;
    input [10:0] input_181;
    input [10:0] input_182;
    input [10:0] input_183;
    input [10:0] input_184;
    input [10:0] input_185;
    input [10:0] input_186;
    input [10:0] input_187;
    input [10:0] input_188;
    input [10:0] input_189;
    input [10:0] input_190;
    input [10:0] input_191;
    input [10:0] input_192;
    input [10:0] input_193;
    input [10:0] input_194;
    input [10:0] input_195;
    input [10:0] input_196;
    input [10:0] input_197;
    input [10:0] input_198;
    input [10:0] input_199;
    input [10:0] input_200;
    input [10:0] input_201;
    input [10:0] input_202;
    input [10:0] input_203;
    input [10:0] input_204;
    input [10:0] input_205;
    input [10:0] input_206;
    input [10:0] input_207;
    input [10:0] input_208;
    input [10:0] input_209;
    input [10:0] input_210;
    input [10:0] input_211;
    input [10:0] input_212;
    input [10:0] input_213;
    input [10:0] input_214;
    input [10:0] input_215;
    input [10:0] input_216;
    input [10:0] input_217;
    input [10:0] input_218;
    input [10:0] input_219;
    input [10:0] input_220;
    input [10:0] input_221;
    input [10:0] input_222;
    input [10:0] input_223;
    input [10:0] input_224;
    input [10:0] input_225;
    input [10:0] input_226;
    input [10:0] input_227;
    input [10:0] input_228;
    input [10:0] input_229;
    input [10:0] input_230;
    input [10:0] input_231;
    input [10:0] input_232;
    input [10:0] input_233;
    input [10:0] input_234;
    input [10:0] input_235;
    input [10:0] input_236;
    input [10:0] input_237;
    input [10:0] input_238;
    input [10:0] input_239;
    input [10:0] input_240;
    input [10:0] input_241;
    input [10:0] input_242;
    input [10:0] input_243;
    input [10:0] input_244;
    input [10:0] input_245;
    input [10:0] input_246;
    input [10:0] input_247;
    input [10:0] input_248;
    input [10:0] input_249;
    input [10:0] input_250;
    input [10:0] input_251;
    input [10:0] input_252;
    input [10:0] input_253;
    input [10:0] input_254;
    input [10:0] input_255;
    input [10:0] input_256;
    input [10:0] input_257;
    input [10:0] input_258;
    input [10:0] input_259;
    input [10:0] input_260;
    input [10:0] input_261;
    input [10:0] input_262;
    input [10:0] input_263;
    input [10:0] input_264;
    input [10:0] input_265;
    input [10:0] input_266;
    input [10:0] input_267;
    input [10:0] input_268;
    input [10:0] input_269;
    input [10:0] input_270;
    input [10:0] input_271;
    input [10:0] input_272;
    input [10:0] input_273;
    input [10:0] input_274;
    input [10:0] input_275;
    input [10:0] input_276;
    input [10:0] input_277;
    input [10:0] input_278;
    input [10:0] input_279;
    input [10:0] input_280;
    input [10:0] input_281;
    input [10:0] input_282;
    input [10:0] input_283;
    input [10:0] input_284;
    input [10:0] input_285;
    input [10:0] input_286;
    input [10:0] input_287;
    input [10:0] input_288;
    input [10:0] input_289;
    input [10:0] input_290;
    input [10:0] input_291;
    input [10:0] input_292;
    input [10:0] input_293;
    input [10:0] input_294;
    input [10:0] input_295;
    input [10:0] input_296;
    input [10:0] input_297;
    input [10:0] input_298;
    input [10:0] input_299;
    input [10:0] input_300;
    input [10:0] input_301;
    input [10:0] input_302;
    input [10:0] input_303;
    input [10:0] input_304;
    input [10:0] input_305;
    input [10:0] input_306;
    input [10:0] input_307;
    input [10:0] input_308;
    input [10:0] input_309;
    input [10:0] input_310;
    input [10:0] input_311;
    input [10:0] input_312;
    input [10:0] input_313;
    input [10:0] input_314;
    input [10:0] input_315;
    input [10:0] input_316;
    input [10:0] input_317;
    input [10:0] input_318;
    input [10:0] input_319;
    input [10:0] input_320;
    input [10:0] input_321;
    input [10:0] input_322;
    input [10:0] input_323;
    input [8:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_v_11_324_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [0:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [44:0] MUX_v_45_2_2;
    input [44:0] input_0;
    input [44:0] input_1;
    input [0:0] sel;
    reg [44:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_45_2_2 = result;
  end
  endfunction


  function automatic [44:0] MUX_v_45_324_2;
    input [44:0] input_0;
    input [44:0] input_1;
    input [44:0] input_2;
    input [44:0] input_3;
    input [44:0] input_4;
    input [44:0] input_5;
    input [44:0] input_6;
    input [44:0] input_7;
    input [44:0] input_8;
    input [44:0] input_9;
    input [44:0] input_10;
    input [44:0] input_11;
    input [44:0] input_12;
    input [44:0] input_13;
    input [44:0] input_14;
    input [44:0] input_15;
    input [44:0] input_16;
    input [44:0] input_17;
    input [44:0] input_18;
    input [44:0] input_19;
    input [44:0] input_20;
    input [44:0] input_21;
    input [44:0] input_22;
    input [44:0] input_23;
    input [44:0] input_24;
    input [44:0] input_25;
    input [44:0] input_26;
    input [44:0] input_27;
    input [44:0] input_28;
    input [44:0] input_29;
    input [44:0] input_30;
    input [44:0] input_31;
    input [44:0] input_32;
    input [44:0] input_33;
    input [44:0] input_34;
    input [44:0] input_35;
    input [44:0] input_36;
    input [44:0] input_37;
    input [44:0] input_38;
    input [44:0] input_39;
    input [44:0] input_40;
    input [44:0] input_41;
    input [44:0] input_42;
    input [44:0] input_43;
    input [44:0] input_44;
    input [44:0] input_45;
    input [44:0] input_46;
    input [44:0] input_47;
    input [44:0] input_48;
    input [44:0] input_49;
    input [44:0] input_50;
    input [44:0] input_51;
    input [44:0] input_52;
    input [44:0] input_53;
    input [44:0] input_54;
    input [44:0] input_55;
    input [44:0] input_56;
    input [44:0] input_57;
    input [44:0] input_58;
    input [44:0] input_59;
    input [44:0] input_60;
    input [44:0] input_61;
    input [44:0] input_62;
    input [44:0] input_63;
    input [44:0] input_64;
    input [44:0] input_65;
    input [44:0] input_66;
    input [44:0] input_67;
    input [44:0] input_68;
    input [44:0] input_69;
    input [44:0] input_70;
    input [44:0] input_71;
    input [44:0] input_72;
    input [44:0] input_73;
    input [44:0] input_74;
    input [44:0] input_75;
    input [44:0] input_76;
    input [44:0] input_77;
    input [44:0] input_78;
    input [44:0] input_79;
    input [44:0] input_80;
    input [44:0] input_81;
    input [44:0] input_82;
    input [44:0] input_83;
    input [44:0] input_84;
    input [44:0] input_85;
    input [44:0] input_86;
    input [44:0] input_87;
    input [44:0] input_88;
    input [44:0] input_89;
    input [44:0] input_90;
    input [44:0] input_91;
    input [44:0] input_92;
    input [44:0] input_93;
    input [44:0] input_94;
    input [44:0] input_95;
    input [44:0] input_96;
    input [44:0] input_97;
    input [44:0] input_98;
    input [44:0] input_99;
    input [44:0] input_100;
    input [44:0] input_101;
    input [44:0] input_102;
    input [44:0] input_103;
    input [44:0] input_104;
    input [44:0] input_105;
    input [44:0] input_106;
    input [44:0] input_107;
    input [44:0] input_108;
    input [44:0] input_109;
    input [44:0] input_110;
    input [44:0] input_111;
    input [44:0] input_112;
    input [44:0] input_113;
    input [44:0] input_114;
    input [44:0] input_115;
    input [44:0] input_116;
    input [44:0] input_117;
    input [44:0] input_118;
    input [44:0] input_119;
    input [44:0] input_120;
    input [44:0] input_121;
    input [44:0] input_122;
    input [44:0] input_123;
    input [44:0] input_124;
    input [44:0] input_125;
    input [44:0] input_126;
    input [44:0] input_127;
    input [44:0] input_128;
    input [44:0] input_129;
    input [44:0] input_130;
    input [44:0] input_131;
    input [44:0] input_132;
    input [44:0] input_133;
    input [44:0] input_134;
    input [44:0] input_135;
    input [44:0] input_136;
    input [44:0] input_137;
    input [44:0] input_138;
    input [44:0] input_139;
    input [44:0] input_140;
    input [44:0] input_141;
    input [44:0] input_142;
    input [44:0] input_143;
    input [44:0] input_144;
    input [44:0] input_145;
    input [44:0] input_146;
    input [44:0] input_147;
    input [44:0] input_148;
    input [44:0] input_149;
    input [44:0] input_150;
    input [44:0] input_151;
    input [44:0] input_152;
    input [44:0] input_153;
    input [44:0] input_154;
    input [44:0] input_155;
    input [44:0] input_156;
    input [44:0] input_157;
    input [44:0] input_158;
    input [44:0] input_159;
    input [44:0] input_160;
    input [44:0] input_161;
    input [44:0] input_162;
    input [44:0] input_163;
    input [44:0] input_164;
    input [44:0] input_165;
    input [44:0] input_166;
    input [44:0] input_167;
    input [44:0] input_168;
    input [44:0] input_169;
    input [44:0] input_170;
    input [44:0] input_171;
    input [44:0] input_172;
    input [44:0] input_173;
    input [44:0] input_174;
    input [44:0] input_175;
    input [44:0] input_176;
    input [44:0] input_177;
    input [44:0] input_178;
    input [44:0] input_179;
    input [44:0] input_180;
    input [44:0] input_181;
    input [44:0] input_182;
    input [44:0] input_183;
    input [44:0] input_184;
    input [44:0] input_185;
    input [44:0] input_186;
    input [44:0] input_187;
    input [44:0] input_188;
    input [44:0] input_189;
    input [44:0] input_190;
    input [44:0] input_191;
    input [44:0] input_192;
    input [44:0] input_193;
    input [44:0] input_194;
    input [44:0] input_195;
    input [44:0] input_196;
    input [44:0] input_197;
    input [44:0] input_198;
    input [44:0] input_199;
    input [44:0] input_200;
    input [44:0] input_201;
    input [44:0] input_202;
    input [44:0] input_203;
    input [44:0] input_204;
    input [44:0] input_205;
    input [44:0] input_206;
    input [44:0] input_207;
    input [44:0] input_208;
    input [44:0] input_209;
    input [44:0] input_210;
    input [44:0] input_211;
    input [44:0] input_212;
    input [44:0] input_213;
    input [44:0] input_214;
    input [44:0] input_215;
    input [44:0] input_216;
    input [44:0] input_217;
    input [44:0] input_218;
    input [44:0] input_219;
    input [44:0] input_220;
    input [44:0] input_221;
    input [44:0] input_222;
    input [44:0] input_223;
    input [44:0] input_224;
    input [44:0] input_225;
    input [44:0] input_226;
    input [44:0] input_227;
    input [44:0] input_228;
    input [44:0] input_229;
    input [44:0] input_230;
    input [44:0] input_231;
    input [44:0] input_232;
    input [44:0] input_233;
    input [44:0] input_234;
    input [44:0] input_235;
    input [44:0] input_236;
    input [44:0] input_237;
    input [44:0] input_238;
    input [44:0] input_239;
    input [44:0] input_240;
    input [44:0] input_241;
    input [44:0] input_242;
    input [44:0] input_243;
    input [44:0] input_244;
    input [44:0] input_245;
    input [44:0] input_246;
    input [44:0] input_247;
    input [44:0] input_248;
    input [44:0] input_249;
    input [44:0] input_250;
    input [44:0] input_251;
    input [44:0] input_252;
    input [44:0] input_253;
    input [44:0] input_254;
    input [44:0] input_255;
    input [44:0] input_256;
    input [44:0] input_257;
    input [44:0] input_258;
    input [44:0] input_259;
    input [44:0] input_260;
    input [44:0] input_261;
    input [44:0] input_262;
    input [44:0] input_263;
    input [44:0] input_264;
    input [44:0] input_265;
    input [44:0] input_266;
    input [44:0] input_267;
    input [44:0] input_268;
    input [44:0] input_269;
    input [44:0] input_270;
    input [44:0] input_271;
    input [44:0] input_272;
    input [44:0] input_273;
    input [44:0] input_274;
    input [44:0] input_275;
    input [44:0] input_276;
    input [44:0] input_277;
    input [44:0] input_278;
    input [44:0] input_279;
    input [44:0] input_280;
    input [44:0] input_281;
    input [44:0] input_282;
    input [44:0] input_283;
    input [44:0] input_284;
    input [44:0] input_285;
    input [44:0] input_286;
    input [44:0] input_287;
    input [44:0] input_288;
    input [44:0] input_289;
    input [44:0] input_290;
    input [44:0] input_291;
    input [44:0] input_292;
    input [44:0] input_293;
    input [44:0] input_294;
    input [44:0] input_295;
    input [44:0] input_296;
    input [44:0] input_297;
    input [44:0] input_298;
    input [44:0] input_299;
    input [44:0] input_300;
    input [44:0] input_301;
    input [44:0] input_302;
    input [44:0] input_303;
    input [44:0] input_304;
    input [44:0] input_305;
    input [44:0] input_306;
    input [44:0] input_307;
    input [44:0] input_308;
    input [44:0] input_309;
    input [44:0] input_310;
    input [44:0] input_311;
    input [44:0] input_312;
    input [44:0] input_313;
    input [44:0] input_314;
    input [44:0] input_315;
    input [44:0] input_316;
    input [44:0] input_317;
    input [44:0] input_318;
    input [44:0] input_319;
    input [44:0] input_320;
    input [44:0] input_321;
    input [44:0] input_322;
    input [44:0] input_323;
    input [8:0] sel;
    reg [44:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_v_45_324_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [54:0] MUX_v_55_2_2;
    input [54:0] input_0;
    input [54:0] input_1;
    input [0:0] sel;
    reg [54:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_55_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] readslicef_10_9_1;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_10_9_1 = tmp[8:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [13:0] signext_14_1;
    input [0:0] vector;
  begin
    signext_14_1= {{13{vector[0]}}, vector};
  end
  endfunction


  function automatic [15:0] signext_16_1;
    input [0:0] vector;
  begin
    signext_16_1= {{15{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input [0:0] vector;
  begin
    signext_5_1= {{4{vector[0]}}, vector};
  end
  endfunction


  function automatic [8:0] signext_9_8;
    input [7:0] vector;
  begin
    signext_9_8= {{1{vector[7]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [57:0] conv_s2s_47_58 ;
    input [46:0]  vector ;
  begin
    conv_s2s_47_58 = {{11{vector[46]}}, vector};
  end
  endfunction


  function automatic [57:0] conv_s2s_57_58 ;
    input [56:0]  vector ;
  begin
    conv_s2s_57_58 = {vector[56], vector};
  end
  endfunction


  function automatic [9:0] conv_s2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_9_17 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_17 = {{8{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [48:0] conv_s2u_47_49 ;
    input [46:0]  vector ;
  begin
    conv_s2u_47_49 = {{2{vector[46]}}, vector};
  end
  endfunction


  function automatic [48:0] conv_s2u_48_49 ;
    input [47:0]  vector ;
  begin
    conv_s2u_48_49 = {vector[47], vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [48:0] conv_u2s_1_49 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_49 = {{48{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_8 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [16:0] conv_u2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_17 =  {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2s_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2s_32_33 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_2_5 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_5 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_3_11 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_11 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_5_13 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_13 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_8_14 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_14 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_11_11 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_11 = vector;
  end
  endfunction


  function automatic [15:0] conv_u2u_11_16 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_16 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_13_13 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_13 = vector;
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction


  function automatic [23:0] conv_u2u_24_24 ;
    input [23:0]  vector ;
  begin
    conv_u2u_24_24 = vector;
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [63:0] conv_u2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_64 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_struct
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_struct (
  clk, rst, conf_info_rsc_dat_batch, conf_info_rsc_dat_n_w, conf_info_rsc_dat_n_h,
      conf_info_rsc_dat_n_c, conf_info_rsc_dat_kern, conf_info_rsc_dat_filt, conf_info_rsc_dat_same,
      conf_info_rsc_dat_stride, conf_info_rsc_vld, conf_info_rsc_rdy, dma_read_ctrl_rsc_dat_size,
      dma_read_ctrl_rsc_dat_length, dma_read_ctrl_rsc_dat_index, dma_read_ctrl_rsc_vld,
      dma_read_ctrl_rsc_rdy, dma_write_ctrl_rsc_dat_size, dma_write_ctrl_rsc_dat_length,
      dma_write_ctrl_rsc_dat_index, dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy,
      dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy, dma_write_chnl_rsc_dat,
      dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, acc_done_rsc_vld
);
  input clk;
  input rst;
  input [31:0] conf_info_rsc_dat_batch;
  input [31:0] conf_info_rsc_dat_n_w;
  input [31:0] conf_info_rsc_dat_n_h;
  input [31:0] conf_info_rsc_dat_n_c;
  input [31:0] conf_info_rsc_dat_kern;
  input [31:0] conf_info_rsc_dat_filt;
  input [31:0] conf_info_rsc_dat_same;
  input [31:0] conf_info_rsc_dat_stride;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [2:0] dma_read_ctrl_rsc_dat_size;
  output [31:0] dma_read_ctrl_rsc_dat_length;
  output [31:0] dma_read_ctrl_rsc_dat_index;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  output [2:0] dma_write_ctrl_rsc_dat_size;
  output [31:0] dma_write_ctrl_rsc_dat_length;
  output [31:0] dma_write_ctrl_rsc_dat_index;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  output acc_done_rsc_vld;


  // Interconnect Declarations
  wire [31:0] plm_in_data_rsci_d_d;
  wire [31:0] plm_in_data_rsci_q_d;
  wire [13:0] plm_in_data_rsci_radr_d;
  wire [13:0] plm_in_data_rsci_wadr_d;
  wire plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_f_data_rsci_d_d;
  wire [31:0] plm_f_data_rsci_q_d;
  wire [15:0] plm_f_data_rsci_radr_d;
  wire [15:0] plm_f_data_rsci_wadr_d;
  wire plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_out_data_rsci_d_d;
  wire [31:0] plm_out_data_rsci_q_d;
  wire [13:0] plm_out_data_rsci_radr_d;
  wire [13:0] plm_out_data_rsci_wadr_d;
  wire plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire plm_in_data_rsc_clken;
  wire [31:0] plm_in_data_rsc_q;
  wire [13:0] plm_in_data_rsc_radr;
  wire plm_in_data_rsc_we;
  wire [31:0] plm_in_data_rsc_d;
  wire [13:0] plm_in_data_rsc_wadr;
  wire plm_f_data_rsc_clken;
  wire [31:0] plm_f_data_rsc_q;
  wire [15:0] plm_f_data_rsc_radr;
  wire plm_f_data_rsc_we;
  wire [31:0] plm_f_data_rsc_d;
  wire [15:0] plm_f_data_rsc_wadr;
  wire plm_out_data_rsc_clken;
  wire [31:0] plm_out_data_rsc_q;
  wire [13:0] plm_out_data_rsc_radr;
  wire plm_out_data_rsc_we;
  wire [31:0] plm_out_data_rsc_d;
  wire [13:0] plm_out_data_rsc_wadr;
  wire [66:0] dma_read_ctrl_rsc_dat;
  wire [66:0] dma_write_ctrl_rsc_dat;
  wire plm_in_data_rsci_we_d_iff;
  wire plm_f_data_rsci_we_d_iff;
  wire plm_out_data_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [255:0] nl_conv2d_cxx_catapult_core_inst_conf_info_rsc_dat;
  assign nl_conv2d_cxx_catapult_core_inst_conf_info_rsc_dat = {conf_info_rsc_dat_batch
      , conf_info_rsc_dat_n_w , conf_info_rsc_dat_n_h , conf_info_rsc_dat_n_c , conf_info_rsc_dat_kern
      , conf_info_rsc_dat_filt , conf_info_rsc_dat_same , conf_info_rsc_dat_stride};
  BLOCK_1R1W_RBW #(.addr_width(32'sd14),
  .data_width(32'sd32),
  .depth(32'sd10368),
  .latency(32'sd1)) plm_in_data_rsc_comp (
      .clk(clk),
      .clken(plm_in_data_rsc_clken),
      .d(plm_in_data_rsc_d),
      .q(plm_in_data_rsc_q),
      .radr(plm_in_data_rsc_radr),
      .wadr(plm_in_data_rsc_wadr),
      .we(plm_in_data_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd16),
  .data_width(32'sd32),
  .depth(32'sd50176),
  .latency(32'sd1)) plm_f_data_rsc_comp (
      .clk(clk),
      .clken(plm_f_data_rsc_clken),
      .d(plm_f_data_rsc_d),
      .q(plm_f_data_rsc_q),
      .radr(plm_f_data_rsc_radr),
      .wadr(plm_f_data_rsc_wadr),
      .we(plm_f_data_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd14),
  .data_width(32'sd32),
  .depth(32'sd10368),
  .latency(32'sd1)) plm_out_data_rsc_comp (
      .clk(clk),
      .clken(plm_out_data_rsc_clken),
      .d(plm_out_data_rsc_d),
      .q(plm_out_data_rsc_q),
      .radr(plm_out_data_rsc_radr),
      .wadr(plm_out_data_rsc_wadr),
      .we(plm_out_data_rsc_we)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_7_14_32_10368_10368_32_1_gen
      plm_in_data_rsci (
      .clken(plm_in_data_rsc_clken),
      .q(plm_in_data_rsc_q),
      .radr(plm_in_data_rsc_radr),
      .we(plm_in_data_rsc_we),
      .d(plm_in_data_rsc_d),
      .wadr(plm_in_data_rsc_wadr),
      .clken_d(1'b1),
      .d_d(plm_in_data_rsci_d_d),
      .q_d(plm_in_data_rsci_q_d),
      .radr_d(plm_in_data_rsci_radr_d),
      .wadr_d(plm_in_data_rsci_wadr_d),
      .we_d(plm_in_data_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_in_data_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_8_16_32_50176_50176_32_1_gen
      plm_f_data_rsci (
      .clken(plm_f_data_rsc_clken),
      .q(plm_f_data_rsc_q),
      .radr(plm_f_data_rsc_radr),
      .we(plm_f_data_rsc_we),
      .d(plm_f_data_rsc_d),
      .wadr(plm_f_data_rsc_wadr),
      .clken_d(1'b1),
      .d_d(plm_f_data_rsci_d_d),
      .q_d(plm_f_data_rsci_q_d),
      .radr_d(plm_f_data_rsci_radr_d),
      .wadr_d(plm_f_data_rsci_wadr_d),
      .we_d(plm_f_data_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_f_data_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_9_14_32_10368_10368_32_1_gen
      plm_out_data_rsci (
      .clken(plm_out_data_rsc_clken),
      .q(plm_out_data_rsc_q),
      .radr(plm_out_data_rsc_radr),
      .we(plm_out_data_rsc_we),
      .d(plm_out_data_rsc_d),
      .wadr(plm_out_data_rsc_wadr),
      .clken_d(1'b1),
      .d_d(plm_out_data_rsci_d_d),
      .q_d(plm_out_data_rsci_q_d),
      .radr_d(plm_out_data_rsci_radr_d),
      .wadr_d(plm_out_data_rsci_wadr_d),
      .we_d(plm_out_data_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_out_data_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core conv2d_cxx_catapult_core_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(nl_conv2d_cxx_catapult_core_inst_conf_info_rsc_dat[255:0]),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .acc_done_rsc_vld(acc_done_rsc_vld),
      .plm_in_data_rsci_d_d(plm_in_data_rsci_d_d),
      .plm_in_data_rsci_q_d(plm_in_data_rsci_q_d),
      .plm_in_data_rsci_radr_d(plm_in_data_rsci_radr_d),
      .plm_in_data_rsci_wadr_d(plm_in_data_rsci_wadr_d),
      .plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_in_data_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_f_data_rsci_d_d(plm_f_data_rsci_d_d),
      .plm_f_data_rsci_q_d(plm_f_data_rsci_q_d),
      .plm_f_data_rsci_radr_d(plm_f_data_rsci_radr_d),
      .plm_f_data_rsci_wadr_d(plm_f_data_rsci_wadr_d),
      .plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_f_data_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_out_data_rsci_d_d(plm_out_data_rsci_d_d),
      .plm_out_data_rsci_q_d(plm_out_data_rsci_q_d),
      .plm_out_data_rsci_radr_d(plm_out_data_rsci_radr_d),
      .plm_out_data_rsci_wadr_d(plm_out_data_rsci_wadr_d),
      .plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_out_data_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_in_data_rsci_we_d_pff(plm_in_data_rsci_we_d_iff),
      .plm_f_data_rsci_we_d_pff(plm_f_data_rsci_we_d_iff),
      .plm_out_data_rsci_we_d_pff(plm_out_data_rsci_we_d_iff)
    );
  assign dma_read_ctrl_rsc_dat_index = dma_read_ctrl_rsc_dat[31:0];
  assign dma_read_ctrl_rsc_dat_length = dma_read_ctrl_rsc_dat[63:32];
  assign dma_read_ctrl_rsc_dat_size = dma_read_ctrl_rsc_dat[66:64];
  assign dma_write_ctrl_rsc_dat_index = dma_write_ctrl_rsc_dat[31:0];
  assign dma_write_ctrl_rsc_dat_length = dma_write_ctrl_rsc_dat[63:32];
  assign dma_write_ctrl_rsc_dat_size = dma_write_ctrl_rsc_dat[66:64];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv2d_cxx_catapult_basic_fx32_dma64
// ------------------------------------------------------------------


module conv2d_cxx_catapult_basic_fx32_dma64 (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, dma_read_ctrl_rsc_dat,
      dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld,
      dma_write_ctrl_rsc_rdy, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy,
      dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, acc_done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  output acc_done_rsc_vld;


  // Interconnect Declarations
  wire [2:0] dma_read_ctrl_rsc_dat_size;
  wire [31:0] dma_read_ctrl_rsc_dat_length;
  wire [31:0] dma_read_ctrl_rsc_dat_index;
  wire [2:0] dma_write_ctrl_rsc_dat_size;
  wire [31:0] dma_write_ctrl_rsc_dat_length;
  wire [31:0] dma_write_ctrl_rsc_dat_index;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_batch;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_batch = conf_info_rsc_dat[255:224];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w = conf_info_rsc_dat[223:192];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h = conf_info_rsc_dat[191:160];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c = conf_info_rsc_dat[159:128];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_kern;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_kern = conf_info_rsc_dat[127:96];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_filt;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_filt = conf_info_rsc_dat[95:64];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_same;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_same = conf_info_rsc_dat[63:32];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_stride;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_stride = conf_info_rsc_dat[31:0];
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_struct conv2d_cxx_catapult_struct_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat_batch(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_batch[31:0]),
      .conf_info_rsc_dat_n_w(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w[31:0]),
      .conf_info_rsc_dat_n_h(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h[31:0]),
      .conf_info_rsc_dat_n_c(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c[31:0]),
      .conf_info_rsc_dat_kern(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_kern[31:0]),
      .conf_info_rsc_dat_filt(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_filt[31:0]),
      .conf_info_rsc_dat_same(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_same[31:0]),
      .conf_info_rsc_dat_stride(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_stride[31:0]),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .dma_read_ctrl_rsc_dat_size(dma_read_ctrl_rsc_dat_size),
      .dma_read_ctrl_rsc_dat_length(dma_read_ctrl_rsc_dat_length),
      .dma_read_ctrl_rsc_dat_index(dma_read_ctrl_rsc_dat_index),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_write_ctrl_rsc_dat_size(dma_write_ctrl_rsc_dat_size),
      .dma_write_ctrl_rsc_dat_length(dma_write_ctrl_rsc_dat_length),
      .dma_write_ctrl_rsc_dat_index(dma_write_ctrl_rsc_dat_index),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .acc_done_rsc_vld(acc_done_rsc_vld)
    );
  assign dma_read_ctrl_rsc_dat = {dma_read_ctrl_rsc_dat_size , dma_read_ctrl_rsc_dat_length
      , dma_read_ctrl_rsc_dat_index};
  assign dma_write_ctrl_rsc_dat = {dma_write_ctrl_rsc_dat_size , dma_write_ctrl_rsc_dat_length
      , dma_write_ctrl_rsc_dat_index};
endmodule



