
//------> ./conv2d_cxx_catapult_ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> ./conv2d_cxx_catapult_ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> ./conv2d_cxx_catapult_ccs_sync_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2d_cxx_catapult_ccs_sync_out_wait_v1 (vld, irdy, ivld, rdy);
  parameter integer rscid = 1;

  input  ivld;
  output irdy;
  output vld;
  input  rdy;

  wire   irdy;
  wire   vld;

  assign vld = ivld;
  assign irdy = rdy;
endmodule

//------> ./conv2d_cxx_catapult_mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./conv2d_cxx_catapult_mgc_in_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_mgc_in_sync_v2 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> ./conv2d_cxx_catapult_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2d_cxx_catapult_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./conv2d_cxx_catapult_ccs_sync_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2d_cxx_catapult_ccs_sync_in_wait_v1 (rdy, vld, irdy, ivld);
  parameter integer rscid = 1;

  output rdy;
  input  vld;
  input  irdy;
  output ivld;

  wire   ivld;
  wire   rdy;

  assign ivld = vld;
  assign rdy = irdy;
endmodule

//------> ./conv2d_cxx_catapult_ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2d_cxx_catapult_ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0

    generate
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> ./conv2d_cxx_catapult_ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module esp_acc_conv2d_cxx_catapult_ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;  // clock enable polarity
    parameter integer ph_arst  = 1;  // async reset polarity
    parameter integer ph_srst  = 1;  // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd;
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
// synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      count = 32'b0;
      peak  = 32'b0;
    end
// synopsys translate_on
  wire din_rdy_drv  ;
  wire dout_vld_drv ;
    wire                 active;
    wire                 din_vld_int;
    wire                 hs_init;

    //assign din_rdy  = din_rdy_drv;    // dout_rdy | (~stat[0] & hs_init);   // original
    assign din_rdy = (fifo_sz > 0) ? (~stat[0] | dout_rdy) && hs_init : dout_rdy ;
    assign dout_vld = dout_vld_drv;
    assign is_idle = (~((din_vld && din_rdy) || (dout_vld && dout_rdy))) && hs_init;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
    assign din_vld_int = din_vld & hs_init;
    assign active =   (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);

      assign din_rdy_drv = dout_rdy | (~stat[0] & hs_init);
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign size_t = (count - {31'b0 , (dout_rdy & stat[fifo_sz-1])}) + { 31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use, no tx)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int  & (~dout_rdy)) // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          if (dout_rdy & stat_behind )
          begin
            // pop n shift
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_nxt & ~((~dout_rdy) & stat[i]))
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0))
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i)%8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]) | ~(active);
          end
        end

        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else
          count_t = n_elem[31:0];
        count = count_t;
// synopsys translate_off
        if ( peak < count )
          peak = count;
// synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      esp_acc_conv2d_cxx_catapult_ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        esp_acc_conv2d_cxx_catapult_ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        esp_acc_conv2d_cxx_catapult_ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
    end
    endgenerate

`ifdef RDY_ASRT
    generate
    if (ph_clk==1)
    begin: POS_CLK_ASSERT

       property rdyAsrt ;
         @(posedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Pos: assert property(rdyAsrt);

    end else if (ph_clk==0)
    begin: NEG_CLK_ASSERT

       property rdyAsrt ;
         @(negedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Neg: assert property(rdyAsrt);

    end
    endgenerate

`endif

endmodule



//------> ./conv2d_cxx_catapult_ccs_pipe_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 */

module esp_acc_conv2d_cxx_catapult_ccs_pipe_v5 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;

// synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = din_vld & !din_rdy;
    assign read_stall  = dout_rdy & !dout_vld;
// synopsys translate_on

    esp_acc_conv2d_cxx_catapult_ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld),
        .din_rdy  (din_rdy),
        .din      (din),
        .dout_vld (dout_vld),
        .dout_rdy (dout_rdy),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ./conv2d_cxx_catapult_ccs_sync_pipe_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_conv2d_cxx_catapult_ccs_sync_pipe_v1 (dout_vld, dout_rdy, din_vld, din_rdy);
  parameter integer rscid = 1;

  input  din_vld;
  output dout_vld;
  input  dout_rdy;
  output din_rdy;

  wire   dout_vld;
  wire   din_rdy;

  assign dout_vld = din_vld;
  assign din_rdy = dout_rdy;
endmodule

//------> /tools/calypto/CATAPULT_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./conv2d_cxx_catapult.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   perenno@esp
//  Generated date: Mon Oct 31 22:33:13 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_cYqiuTts_cns_bctl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_cYqiuTts_cns_bctl (
  clk, rst, plm_outputs_rsc_wadr_ncompute_inst, plm_outputs_rsc_d_ncompute_inst,
      plm_outputs_rsc_we_ncompute_inst, plm_outputs_rsc_req_vz_ncompute_inst, plm_outputs_rsc_we_ncompute_inst_buz,
      conf_info_rsc_rdy_nstore_inst, plm_outputs_rsc_radr_nstore_inst, plm_outputs_rsc_q_nstore_inst,
      plm_outputs_rsc_req_vz_nstore_inst, dma_write_ctrl_rsc_vld_nstore_inst, dma_write_chnl_rsc_vld_nstore_inst,
      done_rsc_vld_nstore_inst, conf_info_rsc_rdy_nstore_inst_bud, plm_outputs_rsc_we_ncompute_inst_buz_bud,
      plm_outputs_rsc_rls_lz_ncompute_inst_bud, plm_outputs_rsc_rls_lz_nstore_inst_bud,
      dma_write_ctrl_rsc_vld_nstore_inst_bud, dma_write_chnl_rsc_vld_nstore_inst_bud,
      done_rsc_vld_nstore_inst_bud, plm_outputs_cns_S0, plm_outputs_cns_R0, plm_outputs_cns_S1,
      plm_outputs_cns_R1, plm_outputs_cns_d_shi0, plm_outputs_cns_d_shi1, plm_outputs_cns_q_sho0,
      plm_outputs_cns_q_sho1, plm_outputs_cns_radr_shi0, plm_outputs_cns_radr_shi1,
      plm_outputs_cns_wadr_shi0, plm_outputs_cns_wadr_shi1, plm_outputs_cns_we_shi0,
      plm_outputs_cns_we_shi1, plm_outputs_rsc_we_ncompute_inst_buz_pff, plm_outputs_rsc_we_ncompute_inst_buz_bud_pff,
      plm_outputs_cns_S0_pff
);
  input clk;
  input rst;
  input [13:0] plm_outputs_rsc_wadr_ncompute_inst;
  input [31:0] plm_outputs_rsc_d_ncompute_inst;
  input plm_outputs_rsc_we_ncompute_inst;
  output plm_outputs_rsc_req_vz_ncompute_inst;
  input plm_outputs_rsc_we_ncompute_inst_buz;
  output conf_info_rsc_rdy_nstore_inst;
  input [13:0] plm_outputs_rsc_radr_nstore_inst;
  output [31:0] plm_outputs_rsc_q_nstore_inst;
  output plm_outputs_rsc_req_vz_nstore_inst;
  output dma_write_ctrl_rsc_vld_nstore_inst;
  output dma_write_chnl_rsc_vld_nstore_inst;
  output done_rsc_vld_nstore_inst;
  input conf_info_rsc_rdy_nstore_inst_bud;
  output plm_outputs_rsc_we_ncompute_inst_buz_bud;
  input plm_outputs_rsc_rls_lz_ncompute_inst_bud;
  input plm_outputs_rsc_rls_lz_nstore_inst_bud;
  input dma_write_ctrl_rsc_vld_nstore_inst_bud;
  input dma_write_chnl_rsc_vld_nstore_inst_bud;
  input done_rsc_vld_nstore_inst_bud;
  output plm_outputs_cns_S0;
  input plm_outputs_cns_R0;
  output plm_outputs_cns_S1;
  input plm_outputs_cns_R1;
  output [31:0] plm_outputs_cns_d_shi0;
  output [31:0] plm_outputs_cns_d_shi1;
  input [31:0] plm_outputs_cns_q_sho0;
  input [31:0] plm_outputs_cns_q_sho1;
  output [13:0] plm_outputs_cns_radr_shi0;
  output [13:0] plm_outputs_cns_radr_shi1;
  output [13:0] plm_outputs_cns_wadr_shi0;
  output [13:0] plm_outputs_cns_wadr_shi1;
  output plm_outputs_cns_we_shi0;
  output plm_outputs_cns_we_shi1;
  input plm_outputs_rsc_we_ncompute_inst_buz_pff;
  output plm_outputs_rsc_we_ncompute_inst_buz_bud_pff;
  output plm_outputs_cns_S0_pff;


  // Interconnect Declarations
  reg plm_outputs_rsc_we_ncompute_inst_buy;
  wire plm_outputs_cns_PC0;
  reg plm_outputs_cns_ppidx;
  reg [1:0] plm_outputs_cns_ppown;
  wire plm_outputs_cns_PC1;
  reg plm_outputs_cns_ppidx_1;
  reg [1:0] plm_outputs_cns_ppown_1;
  wire [1:0] plm_outputs_acc_rmff;
  wire [3:0] nl_plm_outputs_acc_rmff;
  wire plm_outputs_xor_rmff;
  wire [1:0] plm_outputs_acc_1_rmff;
  wire [3:0] nl_plm_outputs_acc_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsc_rdy_nstore_inst = conf_info_rsc_rdy_nstore_inst_bud;
  assign dma_write_ctrl_rsc_vld_nstore_inst = dma_write_ctrl_rsc_vld_nstore_inst_bud;
  assign dma_write_chnl_rsc_vld_nstore_inst = dma_write_chnl_rsc_vld_nstore_inst_bud;
  assign done_rsc_vld_nstore_inst = done_rsc_vld_nstore_inst_bud;
  assign plm_outputs_rsc_req_vz_ncompute_inst = plm_outputs_cns_R0;
  assign plm_outputs_rsc_req_vz_nstore_inst = plm_outputs_cns_R1;
  assign plm_outputs_xor_rmff = plm_outputs_cns_ppidx ^ plm_outputs_cns_PC0;
  assign nl_plm_outputs_acc_rmff = plm_outputs_cns_ppown + conv_u2u_1_2(plm_outputs_cns_PC0)
      + conv_s2u_1_2(plm_outputs_cns_PC1);
  assign plm_outputs_acc_rmff = nl_plm_outputs_acc_rmff[1:0];
  assign plm_outputs_cns_PC0 = plm_outputs_cns_S0 & plm_outputs_rsc_rls_lz_ncompute_inst_bud;
  assign nl_plm_outputs_acc_1_rmff = plm_outputs_cns_ppown_1 + conv_u2u_1_2(plm_outputs_cns_PC1)
      + conv_s2u_1_2(plm_outputs_cns_PC0);
  assign plm_outputs_acc_1_rmff = nl_plm_outputs_acc_1_rmff[1:0];
  assign plm_outputs_cns_PC1 = ((plm_outputs_cns_ppown_1!=2'b00)) & plm_outputs_rsc_rls_lz_nstore_inst_bud;
  assign plm_outputs_rsc_q_nstore_inst = MUX_v_32_2_2(plm_outputs_cns_q_sho0, plm_outputs_cns_q_sho1,
      plm_outputs_cns_ppidx_1);
  assign plm_outputs_cns_d_shi0 = plm_outputs_rsc_d_ncompute_inst;
  assign plm_outputs_cns_radr_shi0 = plm_outputs_rsc_radr_nstore_inst;
  assign plm_outputs_cns_wadr_shi0 = plm_outputs_rsc_wadr_ncompute_inst;
  assign plm_outputs_cns_we_shi0 = plm_outputs_rsc_we_ncompute_inst_buz_pff & plm_outputs_cns_S0_pff
      & (~ plm_outputs_xor_rmff);
  assign plm_outputs_rsc_we_ncompute_inst_buz_bud = plm_outputs_rsc_we_ncompute_inst_buy;
  assign plm_outputs_rsc_we_ncompute_inst_buz_bud_pff = plm_outputs_rsc_we_ncompute_inst;
  assign plm_outputs_cns_S0 = ~((plm_outputs_cns_ppown==2'b10));
  assign plm_outputs_cns_S0_pff = ~((plm_outputs_acc_rmff==2'b10));
  assign plm_outputs_cns_d_shi1 = plm_outputs_rsc_d_ncompute_inst;
  assign plm_outputs_cns_radr_shi1 = plm_outputs_rsc_radr_nstore_inst;
  assign plm_outputs_cns_wadr_shi1 = plm_outputs_rsc_wadr_ncompute_inst;
  assign plm_outputs_cns_we_shi1 = plm_outputs_rsc_we_ncompute_inst_buz_pff & plm_outputs_cns_S0_pff
      & plm_outputs_xor_rmff;
  assign plm_outputs_cns_S1 = (plm_outputs_acc_1_rmff!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsc_we_ncompute_inst_buy <= 1'b0;
      plm_outputs_cns_ppidx <= 1'b0;
      plm_outputs_cns_ppown <= 2'b00;
      plm_outputs_cns_ppidx_1 <= 1'b0;
      plm_outputs_cns_ppown_1 <= 2'b00;
    end
    else begin
      plm_outputs_rsc_we_ncompute_inst_buy <= plm_outputs_rsc_we_ncompute_inst;
      plm_outputs_cns_ppidx <= plm_outputs_xor_rmff;
      plm_outputs_cns_ppown <= plm_outputs_acc_rmff;
      plm_outputs_cns_ppidx_1 <= plm_outputs_cns_ppidx_1 ^ plm_outputs_cns_PC1;
      plm_outputs_cns_ppown_1 <= plm_outputs_acc_1_rmff;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_cYDPQCrs_cns_bctl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_cYDPQCrs_cns_bctl (
  clk, rst, plm_filters_rsc_wadr_nload_inst, plm_filters_rsc_d_nload_inst, plm_filters_rsc_we_nload_inst,
      plm_filters_rsc_req_vz_nload_inst, plm_filters_rsc_we_nload_inst_buz, plm_filters_rsc_radr_ncompute_inst,
      plm_filters_rsc_q_ncompute_inst, plm_filters_rsc_req_vz_ncompute_inst, plm_filters_rsc_we_nload_inst_buz_bud,
      plm_filters_rsc_rls_lz_nload_inst_bud, plm_filters_rsc_rls_lz_ncompute_inst_bud,
      plm_filters_cns_S0, plm_filters_cns_R0, plm_filters_cns_S1, plm_filters_cns_R1,
      plm_filters_cns_d_shi0, plm_filters_cns_d_shi1, plm_filters_cns_q_sho0, plm_filters_cns_q_sho1,
      plm_filters_cns_radr_shi0, plm_filters_cns_radr_shi1, plm_filters_cns_wadr_shi0,
      plm_filters_cns_wadr_shi1, plm_filters_cns_we_shi0, plm_filters_cns_we_shi1,
      plm_filters_rsc_we_nload_inst_buz_pff, plm_filters_rsc_we_nload_inst_buz_bud_pff,
      plm_filters_cns_S0_pff
);
  input clk;
  input rst;
  input [15:0] plm_filters_rsc_wadr_nload_inst;
  input [31:0] plm_filters_rsc_d_nload_inst;
  input plm_filters_rsc_we_nload_inst;
  output plm_filters_rsc_req_vz_nload_inst;
  input plm_filters_rsc_we_nload_inst_buz;
  input [15:0] plm_filters_rsc_radr_ncompute_inst;
  output [31:0] plm_filters_rsc_q_ncompute_inst;
  output plm_filters_rsc_req_vz_ncompute_inst;
  output plm_filters_rsc_we_nload_inst_buz_bud;
  input plm_filters_rsc_rls_lz_nload_inst_bud;
  input plm_filters_rsc_rls_lz_ncompute_inst_bud;
  output plm_filters_cns_S0;
  input plm_filters_cns_R0;
  output plm_filters_cns_S1;
  input plm_filters_cns_R1;
  output [31:0] plm_filters_cns_d_shi0;
  output [31:0] plm_filters_cns_d_shi1;
  input [31:0] plm_filters_cns_q_sho0;
  input [31:0] plm_filters_cns_q_sho1;
  output [15:0] plm_filters_cns_radr_shi0;
  output [15:0] plm_filters_cns_radr_shi1;
  output [15:0] plm_filters_cns_wadr_shi0;
  output [15:0] plm_filters_cns_wadr_shi1;
  output plm_filters_cns_we_shi0;
  output plm_filters_cns_we_shi1;
  input plm_filters_rsc_we_nload_inst_buz_pff;
  output plm_filters_rsc_we_nload_inst_buz_bud_pff;
  output plm_filters_cns_S0_pff;


  // Interconnect Declarations
  reg plm_filters_rsc_we_nload_inst_buy;
  wire plm_filters_cns_PC0;
  reg plm_filters_cns_ppidx;
  reg [1:0] plm_filters_cns_ppown;
  wire plm_filters_cns_PC1;
  reg plm_filters_cns_ppidx_1;
  reg [1:0] plm_filters_cns_ppown_1;
  wire [1:0] plm_filters_acc_rmff;
  wire [3:0] nl_plm_filters_acc_rmff;
  wire plm_filters_xor_rmff;
  wire [1:0] plm_filters_acc_1_rmff;
  wire [3:0] nl_plm_filters_acc_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_req_vz_nload_inst = plm_filters_cns_R0;
  assign plm_filters_rsc_req_vz_ncompute_inst = plm_filters_cns_R1;
  assign plm_filters_xor_rmff = plm_filters_cns_ppidx ^ plm_filters_cns_PC0;
  assign nl_plm_filters_acc_rmff = plm_filters_cns_ppown + conv_u2u_1_2(plm_filters_cns_PC0)
      + conv_s2u_1_2(plm_filters_cns_PC1);
  assign plm_filters_acc_rmff = nl_plm_filters_acc_rmff[1:0];
  assign plm_filters_cns_PC0 = plm_filters_cns_S0 & plm_filters_rsc_rls_lz_nload_inst_bud;
  assign nl_plm_filters_acc_1_rmff = plm_filters_cns_ppown_1 + conv_u2u_1_2(plm_filters_cns_PC1)
      + conv_s2u_1_2(plm_filters_cns_PC0);
  assign plm_filters_acc_1_rmff = nl_plm_filters_acc_1_rmff[1:0];
  assign plm_filters_cns_PC1 = ((plm_filters_cns_ppown_1!=2'b00)) & plm_filters_rsc_rls_lz_ncompute_inst_bud;
  assign plm_filters_rsc_q_ncompute_inst = MUX_v_32_2_2(plm_filters_cns_q_sho0, plm_filters_cns_q_sho1,
      plm_filters_cns_ppidx_1);
  assign plm_filters_cns_d_shi0 = plm_filters_rsc_d_nload_inst;
  assign plm_filters_cns_radr_shi0 = plm_filters_rsc_radr_ncompute_inst;
  assign plm_filters_cns_wadr_shi0 = plm_filters_rsc_wadr_nload_inst;
  assign plm_filters_cns_we_shi0 = plm_filters_rsc_we_nload_inst_buz_pff & plm_filters_cns_S0_pff
      & (~ plm_filters_xor_rmff);
  assign plm_filters_rsc_we_nload_inst_buz_bud = plm_filters_rsc_we_nload_inst_buy;
  assign plm_filters_rsc_we_nload_inst_buz_bud_pff = plm_filters_rsc_we_nload_inst;
  assign plm_filters_cns_S0 = ~((plm_filters_cns_ppown==2'b10));
  assign plm_filters_cns_S0_pff = ~((plm_filters_acc_rmff==2'b10));
  assign plm_filters_cns_d_shi1 = plm_filters_rsc_d_nload_inst;
  assign plm_filters_cns_radr_shi1 = plm_filters_rsc_radr_ncompute_inst;
  assign plm_filters_cns_wadr_shi1 = plm_filters_rsc_wadr_nload_inst;
  assign plm_filters_cns_we_shi1 = plm_filters_rsc_we_nload_inst_buz_pff & plm_filters_cns_S0_pff
      & plm_filters_xor_rmff;
  assign plm_filters_cns_S1 = (plm_filters_acc_1_rmff!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsc_we_nload_inst_buy <= 1'b0;
      plm_filters_cns_ppidx <= 1'b0;
      plm_filters_cns_ppown <= 2'b00;
      plm_filters_cns_ppidx_1 <= 1'b0;
      plm_filters_cns_ppown_1 <= 2'b00;
    end
    else begin
      plm_filters_rsc_we_nload_inst_buy <= plm_filters_rsc_we_nload_inst;
      plm_filters_cns_ppidx <= plm_filters_xor_rmff;
      plm_filters_cns_ppown <= plm_filters_acc_rmff;
      plm_filters_cns_ppidx_1 <= plm_filters_cns_ppidx_1 ^ plm_filters_cns_PC1;
      plm_filters_cns_ppown_1 <= plm_filters_acc_1_rmff;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_cKlrPsts_cns_bctl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_cKlrPsts_cns_bctl (
  clk, rst, conf_info_rsc_rdy_nload_inst, plm_inputs_rsc_wadr_nload_inst, plm_inputs_rsc_d_nload_inst,
      plm_inputs_rsc_we_nload_inst, plm_inputs_rsc_req_vz_nload_inst, dma_read_ctrl_rsc_vld_nload_inst,
      dma_read_chnl_rsc_rdy_nload_inst, done_rsc_vld_nload_inst, plm_filters_rsc_we_nload_inst_buz,
      conf_info_rsc_rdy_ncompute_inst, plm_inputs_rsc_radr_ncompute_inst, plm_inputs_rsc_q_ncompute_inst,
      plm_inputs_rsc_req_vz_ncompute_inst, done_rsc_vld_ncompute_inst, plm_outputs_rsc_we_ncompute_inst_buz,
      conf_info_rsc_rdy_nload_inst_bud, conf_info_rsc_rdy_ncompute_inst_bud, plm_inputs_rsc_rls_lz_nload_inst_bud,
      plm_inputs_rsc_rls_lz_ncompute_inst_bud, plm_filters_rsc_we_nload_inst_buz_bud,
      plm_filters_rsc_rls_lz_nload_inst_bud, plm_filters_rsc_rls_lz_ncompute_inst_bud,
      dma_read_ctrl_rsc_vld_nload_inst_bud, dma_read_chnl_rsc_rdy_nload_inst_bud,
      done_rsc_vld_nload_inst_bud, plm_outputs_rsc_we_ncompute_inst_buz_bud, plm_outputs_rsc_rls_lz_ncompute_inst_bud,
      done_rsc_vld_ncompute_inst_bud, plm_inputs_cns_S0, plm_inputs_cns_R0, plm_inputs_cns_S1,
      plm_inputs_cns_R1, plm_inputs_cns_d_shi0, plm_inputs_cns_d_shi1, plm_inputs_cns_q_sho0,
      plm_inputs_cns_q_sho1, plm_inputs_cns_radr_shi0, plm_inputs_cns_radr_shi1,
      plm_inputs_cns_wadr_shi0, plm_inputs_cns_wadr_shi1, plm_inputs_cns_we_shi0,
      plm_inputs_cns_we_shi1, plm_inputs_cns_S0_pff, plm_filters_rsc_we_nload_inst_buz_pff,
      plm_filters_rsc_we_nload_inst_buz_bud_pff, plm_outputs_rsc_we_ncompute_inst_buz_pff,
      plm_outputs_rsc_we_ncompute_inst_buz_bud_pff
);
  input clk;
  input rst;
  output conf_info_rsc_rdy_nload_inst;
  input [13:0] plm_inputs_rsc_wadr_nload_inst;
  input [31:0] plm_inputs_rsc_d_nload_inst;
  input plm_inputs_rsc_we_nload_inst;
  output plm_inputs_rsc_req_vz_nload_inst;
  output dma_read_ctrl_rsc_vld_nload_inst;
  output dma_read_chnl_rsc_rdy_nload_inst;
  output done_rsc_vld_nload_inst;
  output plm_filters_rsc_we_nload_inst_buz;
  output conf_info_rsc_rdy_ncompute_inst;
  input [13:0] plm_inputs_rsc_radr_ncompute_inst;
  output [31:0] plm_inputs_rsc_q_ncompute_inst;
  output plm_inputs_rsc_req_vz_ncompute_inst;
  output done_rsc_vld_ncompute_inst;
  output plm_outputs_rsc_we_ncompute_inst_buz;
  input conf_info_rsc_rdy_nload_inst_bud;
  input conf_info_rsc_rdy_ncompute_inst_bud;
  input plm_inputs_rsc_rls_lz_nload_inst_bud;
  input plm_inputs_rsc_rls_lz_ncompute_inst_bud;
  input plm_filters_rsc_we_nload_inst_buz_bud;
  input plm_filters_rsc_rls_lz_nload_inst_bud;
  input plm_filters_rsc_rls_lz_ncompute_inst_bud;
  input dma_read_ctrl_rsc_vld_nload_inst_bud;
  input dma_read_chnl_rsc_rdy_nload_inst_bud;
  input done_rsc_vld_nload_inst_bud;
  input plm_outputs_rsc_we_ncompute_inst_buz_bud;
  input plm_outputs_rsc_rls_lz_ncompute_inst_bud;
  input done_rsc_vld_ncompute_inst_bud;
  output plm_inputs_cns_S0;
  input plm_inputs_cns_R0;
  output plm_inputs_cns_S1;
  input plm_inputs_cns_R1;
  output [31:0] plm_inputs_cns_d_shi0;
  output [31:0] plm_inputs_cns_d_shi1;
  input [31:0] plm_inputs_cns_q_sho0;
  input [31:0] plm_inputs_cns_q_sho1;
  output [13:0] plm_inputs_cns_radr_shi0;
  output [13:0] plm_inputs_cns_radr_shi1;
  output [13:0] plm_inputs_cns_wadr_shi0;
  output [13:0] plm_inputs_cns_wadr_shi1;
  output plm_inputs_cns_we_shi0;
  output plm_inputs_cns_we_shi1;
  output plm_inputs_cns_S0_pff;
  output plm_filters_rsc_we_nload_inst_buz_pff;
  input plm_filters_rsc_we_nload_inst_buz_bud_pff;
  output plm_outputs_rsc_we_ncompute_inst_buz_pff;
  input plm_outputs_rsc_we_ncompute_inst_buz_bud_pff;


  // Interconnect Declarations
  wire plm_inputs_cns_PC0;
  reg plm_inputs_cns_ppidx;
  reg [1:0] plm_inputs_cns_ppown;
  wire plm_inputs_cns_PC1;
  reg plm_inputs_cns_ppidx_1;
  reg [1:0] plm_inputs_cns_ppown_1;
  wire [1:0] plm_inputs_acc_rmff;
  wire [3:0] nl_plm_inputs_acc_rmff;
  wire plm_inputs_xor_rmff;
  wire [1:0] plm_inputs_acc_1_rmff;
  wire [3:0] nl_plm_inputs_acc_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsc_rdy_nload_inst = conf_info_rsc_rdy_nload_inst_bud;
  assign conf_info_rsc_rdy_ncompute_inst = conf_info_rsc_rdy_ncompute_inst_bud;
  assign dma_read_ctrl_rsc_vld_nload_inst = dma_read_ctrl_rsc_vld_nload_inst_bud;
  assign dma_read_chnl_rsc_rdy_nload_inst = dma_read_chnl_rsc_rdy_nload_inst_bud;
  assign done_rsc_vld_nload_inst = done_rsc_vld_nload_inst_bud;
  assign done_rsc_vld_ncompute_inst = done_rsc_vld_ncompute_inst_bud;
  assign plm_inputs_rsc_req_vz_nload_inst = plm_inputs_cns_R0;
  assign plm_inputs_rsc_req_vz_ncompute_inst = plm_inputs_cns_R1;
  assign plm_inputs_xor_rmff = plm_inputs_cns_ppidx ^ plm_inputs_cns_PC0;
  assign nl_plm_inputs_acc_rmff = plm_inputs_cns_ppown + conv_u2u_1_2(plm_inputs_cns_PC0)
      + conv_s2u_1_2(plm_inputs_cns_PC1);
  assign plm_inputs_acc_rmff = nl_plm_inputs_acc_rmff[1:0];
  assign plm_inputs_cns_PC0 = plm_inputs_cns_S0 & plm_inputs_rsc_rls_lz_nload_inst_bud;
  assign nl_plm_inputs_acc_1_rmff = plm_inputs_cns_ppown_1 + conv_u2u_1_2(plm_inputs_cns_PC1)
      + conv_s2u_1_2(plm_inputs_cns_PC0);
  assign plm_inputs_acc_1_rmff = nl_plm_inputs_acc_1_rmff[1:0];
  assign plm_inputs_cns_PC1 = ((plm_inputs_cns_ppown_1!=2'b00)) & plm_inputs_rsc_rls_lz_ncompute_inst_bud;
  assign plm_inputs_rsc_q_ncompute_inst = MUX_v_32_2_2(plm_inputs_cns_q_sho0, plm_inputs_cns_q_sho1,
      plm_inputs_cns_ppidx_1);
  assign plm_inputs_cns_d_shi0 = plm_inputs_rsc_d_nload_inst;
  assign plm_inputs_cns_radr_shi0 = plm_inputs_rsc_radr_ncompute_inst;
  assign plm_inputs_cns_wadr_shi0 = plm_inputs_rsc_wadr_nload_inst;
  assign plm_inputs_cns_we_shi0 = plm_inputs_rsc_we_nload_inst & plm_inputs_cns_S0_pff
      & (~ plm_inputs_xor_rmff);
  assign plm_inputs_cns_S0 = ~((plm_inputs_cns_ppown==2'b10));
  assign plm_inputs_cns_S0_pff = ~((plm_inputs_acc_rmff==2'b10));
  assign plm_inputs_cns_d_shi1 = plm_inputs_rsc_d_nload_inst;
  assign plm_inputs_cns_radr_shi1 = plm_inputs_rsc_radr_ncompute_inst;
  assign plm_inputs_cns_wadr_shi1 = plm_inputs_rsc_wadr_nload_inst;
  assign plm_inputs_cns_we_shi1 = plm_inputs_rsc_we_nload_inst & plm_inputs_cns_S0_pff
      & plm_inputs_xor_rmff;
  assign plm_filters_rsc_we_nload_inst_buz = plm_filters_rsc_we_nload_inst_buz_bud;
  assign plm_filters_rsc_we_nload_inst_buz_pff = plm_filters_rsc_we_nload_inst_buz_bud_pff;
  assign plm_outputs_rsc_we_ncompute_inst_buz = plm_outputs_rsc_we_ncompute_inst_buz_bud;
  assign plm_outputs_rsc_we_ncompute_inst_buz_pff = plm_outputs_rsc_we_ncompute_inst_buz_bud_pff;
  assign plm_inputs_cns_S1 = (plm_inputs_acc_1_rmff!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_cns_ppidx <= 1'b0;
      plm_inputs_cns_ppown <= 2'b00;
      plm_inputs_cns_ppidx_1 <= 1'b0;
      plm_inputs_cns_ppown_1 <= 2'b00;
    end
    else begin
      plm_inputs_cns_ppidx <= plm_inputs_xor_rmff;
      plm_inputs_cns_ppown <= plm_inputs_acc_rmff;
      plm_inputs_cns_ppidx_1 <= plm_inputs_cns_ppidx_1 ^ plm_inputs_cns_PC1;
      plm_inputs_cns_ppown_1 <= plm_inputs_acc_1_rmff;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_unreg_hier
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_unreg_hier (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_staller (
  clk, rst, core_wen, core_wten, config_done_cnsi_wen_comp, load_done_cnsi_wen_comp,
      compute_done_cnsi_wen_comp, store_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input config_done_cnsi_wen_comp;
  input load_done_cnsi_wen_comp;
  input compute_done_cnsi_wen_comp;
  input store_done_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = config_done_cnsi_wen_comp & load_done_cnsi_wen_comp & compute_done_cnsi_wen_comp
      & store_done_cnsi_wen_comp;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp
    (
  clk, rst, store_done_cnsi_oswt_unreg, store_done_cnsi_bawt, store_done_cnsi_wen_comp,
      store_done_cnsi_biwt, store_done_cnsi_bdwt, store_done_cnsi_bcwt
);
  input clk;
  input rst;
  input store_done_cnsi_oswt_unreg;
  output store_done_cnsi_bawt;
  output store_done_cnsi_wen_comp;
  input store_done_cnsi_biwt;
  input store_done_cnsi_bdwt;
  output store_done_cnsi_bcwt;
  reg store_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign store_done_cnsi_bawt = store_done_cnsi_biwt | store_done_cnsi_bcwt;
  assign store_done_cnsi_wen_comp = (~ store_done_cnsi_oswt_unreg) | store_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      store_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      store_done_cnsi_bcwt <= ~((~(store_done_cnsi_bcwt | store_done_cnsi_biwt))
          | store_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl
    (
  core_wen, store_done_cnsi_oswt_unreg, store_done_cnsi_iswt0, store_done_cnsi_ivld,
      store_done_cnsi_biwt, store_done_cnsi_bdwt, store_done_cnsi_bcwt, store_done_cnsi_irdy_core_sct
);
  input core_wen;
  input store_done_cnsi_oswt_unreg;
  input store_done_cnsi_iswt0;
  input store_done_cnsi_ivld;
  output store_done_cnsi_biwt;
  output store_done_cnsi_bdwt;
  input store_done_cnsi_bcwt;
  output store_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire store_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign store_done_cnsi_bdwt = store_done_cnsi_oswt_unreg & core_wen;
  assign store_done_cnsi_biwt = store_done_cnsi_ogwt & store_done_cnsi_ivld;
  assign store_done_cnsi_ogwt = store_done_cnsi_iswt0 & (~ store_done_cnsi_bcwt);
  assign store_done_cnsi_irdy_core_sct = store_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp
    (
  clk, rst, compute_done_cnsi_oswt_unreg, compute_done_cnsi_bawt, compute_done_cnsi_wen_comp,
      compute_done_cnsi_biwt, compute_done_cnsi_bdwt, compute_done_cnsi_bcwt
);
  input clk;
  input rst;
  input compute_done_cnsi_oswt_unreg;
  output compute_done_cnsi_bawt;
  output compute_done_cnsi_wen_comp;
  input compute_done_cnsi_biwt;
  input compute_done_cnsi_bdwt;
  output compute_done_cnsi_bcwt;
  reg compute_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign compute_done_cnsi_bawt = compute_done_cnsi_biwt | compute_done_cnsi_bcwt;
  assign compute_done_cnsi_wen_comp = (~ compute_done_cnsi_oswt_unreg) | compute_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      compute_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      compute_done_cnsi_bcwt <= ~((~(compute_done_cnsi_bcwt | compute_done_cnsi_biwt))
          | compute_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl
    (
  core_wen, compute_done_cnsi_oswt_unreg, compute_done_cnsi_iswt0, compute_done_cnsi_ivld,
      compute_done_cnsi_biwt, compute_done_cnsi_bdwt, compute_done_cnsi_bcwt, compute_done_cnsi_irdy_core_sct
);
  input core_wen;
  input compute_done_cnsi_oswt_unreg;
  input compute_done_cnsi_iswt0;
  input compute_done_cnsi_ivld;
  output compute_done_cnsi_biwt;
  output compute_done_cnsi_bdwt;
  input compute_done_cnsi_bcwt;
  output compute_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire compute_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign compute_done_cnsi_bdwt = compute_done_cnsi_oswt_unreg & core_wen;
  assign compute_done_cnsi_biwt = compute_done_cnsi_ogwt & compute_done_cnsi_ivld;
  assign compute_done_cnsi_ogwt = compute_done_cnsi_iswt0 & (~ compute_done_cnsi_bcwt);
  assign compute_done_cnsi_irdy_core_sct = compute_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp
    (
  clk, rst, load_done_cnsi_oswt_unreg, load_done_cnsi_bawt, load_done_cnsi_wen_comp,
      load_done_cnsi_biwt, load_done_cnsi_bdwt, load_done_cnsi_bcwt
);
  input clk;
  input rst;
  input load_done_cnsi_oswt_unreg;
  output load_done_cnsi_bawt;
  output load_done_cnsi_wen_comp;
  input load_done_cnsi_biwt;
  input load_done_cnsi_bdwt;
  output load_done_cnsi_bcwt;
  reg load_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign load_done_cnsi_bawt = load_done_cnsi_biwt | load_done_cnsi_bcwt;
  assign load_done_cnsi_wen_comp = (~ load_done_cnsi_oswt_unreg) | load_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      load_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      load_done_cnsi_bcwt <= ~((~(load_done_cnsi_bcwt | load_done_cnsi_biwt)) | load_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl
    (
  core_wen, load_done_cnsi_oswt_unreg, load_done_cnsi_iswt0, load_done_cnsi_irdy_core_psct,
      load_done_cnsi_ivld, load_done_cnsi_biwt, load_done_cnsi_bdwt, load_done_cnsi_bcwt,
      load_done_cnsi_irdy_core_sct
);
  input core_wen;
  input load_done_cnsi_oswt_unreg;
  input load_done_cnsi_iswt0;
  input load_done_cnsi_irdy_core_psct;
  input load_done_cnsi_ivld;
  output load_done_cnsi_biwt;
  output load_done_cnsi_bdwt;
  input load_done_cnsi_bcwt;
  output load_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire load_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign load_done_cnsi_bdwt = load_done_cnsi_oswt_unreg & core_wen;
  assign load_done_cnsi_biwt = load_done_cnsi_ogwt & load_done_cnsi_ivld;
  assign load_done_cnsi_ogwt = load_done_cnsi_iswt0 & (~ load_done_cnsi_bcwt);
  assign load_done_cnsi_irdy_core_sct = load_done_cnsi_irdy_core_psct & load_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp
    (
  clk, rst, config_done_cnsi_oswt_unreg, config_done_cnsi_bawt, config_done_cnsi_wen_comp,
      config_done_cnsi_biwt, config_done_cnsi_bdwt, config_done_cnsi_bcwt
);
  input clk;
  input rst;
  input config_done_cnsi_oswt_unreg;
  output config_done_cnsi_bawt;
  output config_done_cnsi_wen_comp;
  input config_done_cnsi_biwt;
  input config_done_cnsi_bdwt;
  output config_done_cnsi_bcwt;
  reg config_done_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign config_done_cnsi_bawt = config_done_cnsi_biwt | config_done_cnsi_bcwt;
  assign config_done_cnsi_wen_comp = (~ config_done_cnsi_oswt_unreg) | config_done_cnsi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      config_done_cnsi_bcwt <= 1'b0;
    end
    else begin
      config_done_cnsi_bcwt <= ~((~(config_done_cnsi_bcwt | config_done_cnsi_biwt))
          | config_done_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl
    (
  core_wen, config_done_cnsi_oswt_unreg, config_done_cnsi_iswt0, config_done_cnsi_ivld,
      config_done_cnsi_biwt, config_done_cnsi_bdwt, config_done_cnsi_bcwt, config_done_cnsi_irdy_core_sct
);
  input core_wen;
  input config_done_cnsi_oswt_unreg;
  input config_done_cnsi_iswt0;
  input config_done_cnsi_ivld;
  output config_done_cnsi_biwt;
  output config_done_cnsi_bdwt;
  input config_done_cnsi_bcwt;
  output config_done_cnsi_irdy_core_sct;


  // Interconnect Declarations
  wire config_done_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign config_done_cnsi_bdwt = config_done_cnsi_oswt_unreg & core_wen;
  assign config_done_cnsi_biwt = config_done_cnsi_ogwt & config_done_cnsi_ivld;
  assign config_done_cnsi_ogwt = config_done_cnsi_iswt0 & (~ config_done_cnsi_bcwt);
  assign config_done_cnsi_irdy_core_sct = config_done_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp
    (
  clk, rst, acc_done_rsci_bawt, acc_done_rsci_biwt, acc_done_rsci_bdwt
);
  input clk;
  input rst;
  output acc_done_rsci_bawt;
  input acc_done_rsci_biwt;
  input acc_done_rsci_bdwt;


  // Interconnect Declarations
  reg acc_done_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign acc_done_rsci_bawt = acc_done_rsci_biwt | acc_done_rsci_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      acc_done_rsci_bcwt <= 1'b0;
    end
    else begin
      acc_done_rsci_bcwt <= ~((~(acc_done_rsci_bcwt | acc_done_rsci_biwt)) | acc_done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl
    (
  core_wen, acc_done_rsci_oswt_unreg, acc_done_rsci_iswt0, core_wten, acc_done_rsci_biwt,
      acc_done_rsci_bdwt
);
  input core_wen;
  input acc_done_rsci_oswt_unreg;
  input acc_done_rsci_iswt0;
  input core_wten;
  output acc_done_rsci_biwt;
  output acc_done_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign acc_done_rsci_bdwt = acc_done_rsci_oswt_unreg & core_wen;
  assign acc_done_rsci_biwt = (~ core_wten) & acc_done_rsci_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2d_cxx_catapult_config_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2d_cxx_catapult_config_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_staller (
  core_wen, conf_info_rsci_wen_comp, plm_conf_load_rsci_wen_comp, plm_conf_compute_rsci_wen_comp,
      plm_conf_store_rsci_wen_comp, done_rsci_wen_comp
);
  output core_wen;
  input conf_info_rsci_wen_comp;
  input plm_conf_load_rsci_wen_comp;
  input plm_conf_compute_rsci_wen_comp;
  input plm_conf_store_rsci_wen_comp;
  input done_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & plm_conf_load_rsci_wen_comp & plm_conf_compute_rsci_wen_comp
      & plm_conf_store_rsci_wen_comp & done_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt_unreg, done_rsci_bawt, done_rsci_wen_comp, done_rsci_biwt,
      done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bawt = done_rsci_biwt | done_rsci_bcwt;
  assign done_rsci_wen_comp = (~ done_rsci_oswt_unreg) | done_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt_unreg, done_rsci_iswt0, done_rsci_biwt, done_rsci_bdwt,
      done_rsci_bcwt, done_rsci_ivld_core_sct, done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt_unreg;
  input done_rsci_iswt0;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt_unreg & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_iswt0 & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_dp
    (
  clk, rst, plm_conf_store_rsci_oswt_unreg, plm_conf_store_rsci_bawt, plm_conf_store_rsci_wen_comp,
      plm_conf_store_rsci_biwt, plm_conf_store_rsci_bdwt, plm_conf_store_rsci_bcwt
);
  input clk;
  input rst;
  input plm_conf_store_rsci_oswt_unreg;
  output plm_conf_store_rsci_bawt;
  output plm_conf_store_rsci_wen_comp;
  input plm_conf_store_rsci_biwt;
  input plm_conf_store_rsci_bdwt;
  output plm_conf_store_rsci_bcwt;
  reg plm_conf_store_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_store_rsci_bawt = plm_conf_store_rsci_biwt | plm_conf_store_rsci_bcwt;
  assign plm_conf_store_rsci_wen_comp = (~ plm_conf_store_rsci_oswt_unreg) | plm_conf_store_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_store_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_conf_store_rsci_bcwt <= ~((~(plm_conf_store_rsci_bcwt | plm_conf_store_rsci_biwt))
          | plm_conf_store_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl
    (
  core_wen, plm_conf_store_rsci_oswt_unreg, plm_conf_store_rsci_iswt0, plm_conf_store_rsci_irdy,
      plm_conf_store_rsci_biwt, plm_conf_store_rsci_bdwt, plm_conf_store_rsci_bcwt,
      plm_conf_store_rsci_ivld_core_sct
);
  input core_wen;
  input plm_conf_store_rsci_oswt_unreg;
  input plm_conf_store_rsci_iswt0;
  input plm_conf_store_rsci_irdy;
  output plm_conf_store_rsci_biwt;
  output plm_conf_store_rsci_bdwt;
  input plm_conf_store_rsci_bcwt;
  output plm_conf_store_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire plm_conf_store_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_store_rsci_bdwt = plm_conf_store_rsci_oswt_unreg & core_wen;
  assign plm_conf_store_rsci_biwt = plm_conf_store_rsci_ogwt & plm_conf_store_rsci_irdy;
  assign plm_conf_store_rsci_ogwt = plm_conf_store_rsci_iswt0 & (~ plm_conf_store_rsci_bcwt);
  assign plm_conf_store_rsci_ivld_core_sct = plm_conf_store_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp
    (
  clk, rst, plm_conf_compute_rsci_oswt_unreg, plm_conf_compute_rsci_bawt, plm_conf_compute_rsci_wen_comp,
      plm_conf_compute_rsci_biwt, plm_conf_compute_rsci_bdwt, plm_conf_compute_rsci_bcwt
);
  input clk;
  input rst;
  input plm_conf_compute_rsci_oswt_unreg;
  output plm_conf_compute_rsci_bawt;
  output plm_conf_compute_rsci_wen_comp;
  input plm_conf_compute_rsci_biwt;
  input plm_conf_compute_rsci_bdwt;
  output plm_conf_compute_rsci_bcwt;
  reg plm_conf_compute_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_compute_rsci_bawt = plm_conf_compute_rsci_biwt | plm_conf_compute_rsci_bcwt;
  assign plm_conf_compute_rsci_wen_comp = (~ plm_conf_compute_rsci_oswt_unreg) |
      plm_conf_compute_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_compute_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_conf_compute_rsci_bcwt <= ~((~(plm_conf_compute_rsci_bcwt | plm_conf_compute_rsci_biwt))
          | plm_conf_compute_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl
    (
  core_wen, plm_conf_compute_rsci_oswt_unreg, plm_conf_compute_rsci_iswt0, plm_conf_compute_rsci_irdy,
      plm_conf_compute_rsci_biwt, plm_conf_compute_rsci_bdwt, plm_conf_compute_rsci_bcwt,
      plm_conf_compute_rsci_ivld_core_sct
);
  input core_wen;
  input plm_conf_compute_rsci_oswt_unreg;
  input plm_conf_compute_rsci_iswt0;
  input plm_conf_compute_rsci_irdy;
  output plm_conf_compute_rsci_biwt;
  output plm_conf_compute_rsci_bdwt;
  input plm_conf_compute_rsci_bcwt;
  output plm_conf_compute_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire plm_conf_compute_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_compute_rsci_bdwt = plm_conf_compute_rsci_oswt_unreg & core_wen;
  assign plm_conf_compute_rsci_biwt = plm_conf_compute_rsci_ogwt & plm_conf_compute_rsci_irdy;
  assign plm_conf_compute_rsci_ogwt = plm_conf_compute_rsci_iswt0 & (~ plm_conf_compute_rsci_bcwt);
  assign plm_conf_compute_rsci_ivld_core_sct = plm_conf_compute_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_dp
    (
  clk, rst, plm_conf_load_rsci_oswt_unreg, plm_conf_load_rsci_bawt, plm_conf_load_rsci_wen_comp,
      plm_conf_load_rsci_biwt, plm_conf_load_rsci_bdwt, plm_conf_load_rsci_bcwt
);
  input clk;
  input rst;
  input plm_conf_load_rsci_oswt_unreg;
  output plm_conf_load_rsci_bawt;
  output plm_conf_load_rsci_wen_comp;
  input plm_conf_load_rsci_biwt;
  input plm_conf_load_rsci_bdwt;
  output plm_conf_load_rsci_bcwt;
  reg plm_conf_load_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_load_rsci_bawt = plm_conf_load_rsci_biwt | plm_conf_load_rsci_bcwt;
  assign plm_conf_load_rsci_wen_comp = (~ plm_conf_load_rsci_oswt_unreg) | plm_conf_load_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_load_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_conf_load_rsci_bcwt <= ~((~(plm_conf_load_rsci_bcwt | plm_conf_load_rsci_biwt))
          | plm_conf_load_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl
    (
  core_wen, plm_conf_load_rsci_oswt_unreg, plm_conf_load_rsci_iswt0, plm_conf_load_rsci_irdy,
      plm_conf_load_rsci_biwt, plm_conf_load_rsci_bdwt, plm_conf_load_rsci_bcwt,
      plm_conf_load_rsci_ivld_core_sct
);
  input core_wen;
  input plm_conf_load_rsci_oswt_unreg;
  input plm_conf_load_rsci_iswt0;
  input plm_conf_load_rsci_irdy;
  output plm_conf_load_rsci_biwt;
  output plm_conf_load_rsci_bdwt;
  input plm_conf_load_rsci_bcwt;
  output plm_conf_load_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire plm_conf_load_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_conf_load_rsci_bdwt = plm_conf_load_rsci_oswt_unreg & core_wen;
  assign plm_conf_load_rsci_biwt = plm_conf_load_rsci_ogwt & plm_conf_load_rsci_irdy;
  assign plm_conf_load_rsci_ogwt = plm_conf_load_rsci_iswt0 & (~ plm_conf_load_rsci_bcwt);
  assign plm_conf_load_rsci_ivld_core_sct = plm_conf_load_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_dp (
  clk, rst, conf_info_rsci_oswt_unreg, conf_info_rsci_bawt, conf_info_rsci_wen_comp,
      conf_info_rsci_idat_mxwt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  output conf_info_rsci_wen_comp;
  output [255:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  reg [255:0] conf_info_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bawt = conf_info_rsci_biwt | conf_info_rsci_bcwt;
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt_unreg) | conf_info_rsci_bawt;
  assign conf_info_rsci_idat_mxwt = MUX_v_256_2_2(conf_info_rsci_idat, conf_info_rsci_idat_bfwt,
      conf_info_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt <= conf_info_rsci_idat;
    end
  end

  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt_unreg, conf_info_rsci_iswt0, conf_info_rsci_biwt,
      conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt_unreg & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_iswt0 & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_8_16_32_50176_50176_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_8_16_32_50176_50176_32_1_gen
    (
  we, d, wadr, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [31:0] d;
  output [15:0] wadr;
  input [31:0] d_d;
  input [15:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_7_14_32_10368_10368_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_7_14_32_10368_10368_32_1_gen
    (
  we, d, wadr, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2d_cxx_catapult_load_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2d_cxx_catapult_load_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_staller (
  clk, rst, core_wen, core_wten, conf_info_rsci_wen_comp, dma_read_chnl_rsci_wen_comp,
      done_rsci_wen_comp, plm_inputs_rsc_req_obj_wen_comp, plm_filters_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input conf_info_rsci_wen_comp;
  input dma_read_chnl_rsci_wen_comp;
  input done_rsci_wen_comp;
  input plm_inputs_rsc_req_obj_wen_comp;
  input plm_filters_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & dma_read_chnl_rsci_wen_comp & done_rsci_wen_comp
      & plm_inputs_rsc_req_obj_wen_comp & plm_filters_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp
    (
  clk, rst, plm_filters_rsc_req_obj_oswt_unreg, plm_filters_rsc_req_obj_bawt, plm_filters_rsc_req_obj_wen_comp,
      plm_filters_rsc_req_obj_biwt, plm_filters_rsc_req_obj_bdwt, plm_filters_rsc_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_filters_rsc_req_obj_oswt_unreg;
  output plm_filters_rsc_req_obj_bawt;
  output plm_filters_rsc_req_obj_wen_comp;
  input plm_filters_rsc_req_obj_biwt;
  input plm_filters_rsc_req_obj_bdwt;
  output plm_filters_rsc_req_obj_bcwt;
  reg plm_filters_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_req_obj_bawt = plm_filters_rsc_req_obj_biwt | plm_filters_rsc_req_obj_bcwt;
  assign plm_filters_rsc_req_obj_wen_comp = (~ plm_filters_rsc_req_obj_oswt_unreg)
      | plm_filters_rsc_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_filters_rsc_req_obj_bcwt <= ~((~(plm_filters_rsc_req_obj_bcwt | plm_filters_rsc_req_obj_biwt))
          | plm_filters_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl
    (
  core_wen, plm_filters_rsc_req_obj_oswt_unreg, plm_filters_rsc_req_obj_iswt0, plm_filters_rsc_req_obj_vd,
      plm_filters_rsc_req_obj_biwt, plm_filters_rsc_req_obj_bdwt, plm_filters_rsc_req_obj_bcwt
);
  input core_wen;
  input plm_filters_rsc_req_obj_oswt_unreg;
  input plm_filters_rsc_req_obj_iswt0;
  input plm_filters_rsc_req_obj_vd;
  output plm_filters_rsc_req_obj_biwt;
  output plm_filters_rsc_req_obj_bdwt;
  input plm_filters_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_req_obj_bdwt = plm_filters_rsc_req_obj_oswt_unreg & core_wen;
  assign plm_filters_rsc_req_obj_biwt = plm_filters_rsc_req_obj_iswt0 & (~ plm_filters_rsc_req_obj_bcwt)
      & plm_filters_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp
    (
  clk, rst, plm_inputs_rsc_req_obj_oswt_unreg, plm_inputs_rsc_req_obj_bawt, plm_inputs_rsc_req_obj_wen_comp,
      plm_inputs_rsc_req_obj_biwt, plm_inputs_rsc_req_obj_bdwt, plm_inputs_rsc_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_inputs_rsc_req_obj_oswt_unreg;
  output plm_inputs_rsc_req_obj_bawt;
  output plm_inputs_rsc_req_obj_wen_comp;
  input plm_inputs_rsc_req_obj_biwt;
  input plm_inputs_rsc_req_obj_bdwt;
  output plm_inputs_rsc_req_obj_bcwt;
  reg plm_inputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_req_obj_bawt = plm_inputs_rsc_req_obj_biwt | plm_inputs_rsc_req_obj_bcwt;
  assign plm_inputs_rsc_req_obj_wen_comp = (~ plm_inputs_rsc_req_obj_oswt_unreg)
      | plm_inputs_rsc_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_inputs_rsc_req_obj_bcwt <= ~((~(plm_inputs_rsc_req_obj_bcwt | plm_inputs_rsc_req_obj_biwt))
          | plm_inputs_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl
    (
  core_wen, plm_inputs_rsc_req_obj_oswt_unreg, plm_inputs_rsc_req_obj_iswt0, plm_inputs_rsc_req_obj_vd,
      plm_inputs_rsc_req_obj_biwt, plm_inputs_rsc_req_obj_bdwt, plm_inputs_rsc_req_obj_bcwt
);
  input core_wen;
  input plm_inputs_rsc_req_obj_oswt_unreg;
  input plm_inputs_rsc_req_obj_iswt0;
  input plm_inputs_rsc_req_obj_vd;
  output plm_inputs_rsc_req_obj_biwt;
  output plm_inputs_rsc_req_obj_bdwt;
  input plm_inputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_req_obj_bdwt = plm_inputs_rsc_req_obj_oswt_unreg & core_wen;
  assign plm_inputs_rsc_req_obj_biwt = plm_inputs_rsc_req_obj_iswt0 & (~ plm_inputs_rsc_req_obj_bcwt)
      & plm_inputs_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp
    (
  clk, rst, plm_filters_rsc_rls_obj_bawt, plm_filters_rsc_rls_obj_biwt, plm_filters_rsc_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_filters_rsc_rls_obj_bawt;
  input plm_filters_rsc_rls_obj_biwt;
  input plm_filters_rsc_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_filters_rsc_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_rls_obj_bawt = plm_filters_rsc_rls_obj_biwt | plm_filters_rsc_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsc_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_filters_rsc_rls_obj_bcwt <= ~((~(plm_filters_rsc_rls_obj_bcwt | plm_filters_rsc_rls_obj_biwt))
          | plm_filters_rsc_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl
    (
  core_wen, core_wten, plm_filters_rsc_rls_obj_oswt_unreg, plm_filters_rsc_rls_obj_iswt0,
      plm_filters_rsc_rls_obj_biwt, plm_filters_rsc_rls_obj_bdwt
);
  input core_wen;
  input core_wten;
  input plm_filters_rsc_rls_obj_oswt_unreg;
  input plm_filters_rsc_rls_obj_iswt0;
  output plm_filters_rsc_rls_obj_biwt;
  output plm_filters_rsc_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_rls_obj_bdwt = plm_filters_rsc_rls_obj_oswt_unreg & core_wen;
  assign plm_filters_rsc_rls_obj_biwt = (~ core_wten) & plm_filters_rsc_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp
    (
  clk, rst, plm_inputs_rsc_rls_obj_bawt, plm_inputs_rsc_rls_obj_biwt, plm_inputs_rsc_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_inputs_rsc_rls_obj_bawt;
  input plm_inputs_rsc_rls_obj_biwt;
  input plm_inputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_inputs_rsc_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_rls_obj_bawt = plm_inputs_rsc_rls_obj_biwt | plm_inputs_rsc_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsc_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_inputs_rsc_rls_obj_bcwt <= ~((~(plm_inputs_rsc_rls_obj_bcwt | plm_inputs_rsc_rls_obj_biwt))
          | plm_inputs_rsc_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl
    (
  core_wen, core_wten, plm_inputs_rsc_rls_obj_oswt_unreg, plm_inputs_rsc_rls_obj_iswt0,
      plm_inputs_rsc_rls_obj_biwt, plm_inputs_rsc_rls_obj_bdwt
);
  input core_wen;
  input core_wten;
  input plm_inputs_rsc_rls_obj_oswt_unreg;
  input plm_inputs_rsc_rls_obj_iswt0;
  output plm_inputs_rsc_rls_obj_biwt;
  output plm_inputs_rsc_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_rls_obj_bdwt = plm_inputs_rsc_rls_obj_oswt_unreg & core_wen;
  assign plm_inputs_rsc_rls_obj_biwt = (~ core_wten) & plm_inputs_rsc_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt_unreg, done_rsci_bawt, done_rsci_wen_comp, done_rsci_biwt,
      done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bawt = done_rsci_biwt | done_rsci_bcwt;
  assign done_rsci_wen_comp = (~ done_rsci_oswt_unreg) | done_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt_unreg, done_rsci_iswt0, done_rsci_biwt, done_rsci_bdwt,
      done_rsci_bcwt, done_rsci_ivld_core_sct, done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt_unreg;
  input done_rsci_iswt0;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt_unreg & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_iswt0 & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
    (
  clk, rst, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_bawt, dma_read_chnl_rsci_wen_comp,
      dma_read_chnl_rsci_idat_mxwt, dma_read_chnl_rsci_biwt, dma_read_chnl_rsci_bdwt,
      dma_read_chnl_rsci_bcwt, dma_read_chnl_rsci_idat
);
  input clk;
  input rst;
  input dma_read_chnl_rsci_oswt_unreg;
  output dma_read_chnl_rsci_bawt;
  output dma_read_chnl_rsci_wen_comp;
  output [31:0] dma_read_chnl_rsci_idat_mxwt;
  input dma_read_chnl_rsci_biwt;
  input dma_read_chnl_rsci_bdwt;
  output dma_read_chnl_rsci_bcwt;
  reg dma_read_chnl_rsci_bcwt;
  input [63:0] dma_read_chnl_rsci_idat;


  // Interconnect Declarations
  reg [31:0] dma_read_chnl_rsci_idat_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_rsci_bawt = dma_read_chnl_rsci_biwt | dma_read_chnl_rsci_bcwt;
  assign dma_read_chnl_rsci_wen_comp = (~ dma_read_chnl_rsci_oswt_unreg) | dma_read_chnl_rsci_bawt;
  assign dma_read_chnl_rsci_idat_mxwt = MUX_v_32_2_2((dma_read_chnl_rsci_idat[31:0]),
      dma_read_chnl_rsci_idat_bfwt_31_0, dma_read_chnl_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_read_chnl_rsci_bcwt <= ~((~(dma_read_chnl_rsci_bcwt | dma_read_chnl_rsci_biwt))
          | dma_read_chnl_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_rsci_idat_bfwt_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( dma_read_chnl_rsci_biwt ) begin
      dma_read_chnl_rsci_idat_bfwt_31_0 <= dma_read_chnl_rsci_idat[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
    (
  core_wen, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_iswt0, dma_read_chnl_rsci_biwt,
      dma_read_chnl_rsci_bdwt, dma_read_chnl_rsci_bcwt, dma_read_chnl_rsci_irdy_core_sct,
      dma_read_chnl_rsci_ivld
);
  input core_wen;
  input dma_read_chnl_rsci_oswt_unreg;
  input dma_read_chnl_rsci_iswt0;
  output dma_read_chnl_rsci_biwt;
  output dma_read_chnl_rsci_bdwt;
  input dma_read_chnl_rsci_bcwt;
  output dma_read_chnl_rsci_irdy_core_sct;
  input dma_read_chnl_rsci_ivld;


  // Interconnect Declarations
  wire dma_read_chnl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_rsci_bdwt = dma_read_chnl_rsci_oswt_unreg & core_wen;
  assign dma_read_chnl_rsci_biwt = dma_read_chnl_rsci_ogwt & dma_read_chnl_rsci_ivld;
  assign dma_read_chnl_rsci_ogwt = dma_read_chnl_rsci_iswt0 & (~ dma_read_chnl_rsci_bcwt);
  assign dma_read_chnl_rsci_irdy_core_sct = dma_read_chnl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
    (
  clk, rst, dma_read_ctrl_rsci_bawt, dma_read_ctrl_rsci_irdy_mxwt, dma_read_ctrl_rsci_irdy,
      dma_read_ctrl_rsci_biwt, dma_read_ctrl_rsci_bdwt
);
  input clk;
  input rst;
  output dma_read_ctrl_rsci_bawt;
  output dma_read_ctrl_rsci_irdy_mxwt;
  input dma_read_ctrl_rsci_irdy;
  input dma_read_ctrl_rsci_biwt;
  input dma_read_ctrl_rsci_bdwt;


  // Interconnect Declarations
  reg dma_read_ctrl_rsci_bcwt;
  reg dma_read_ctrl_rsci_irdy_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_rsci_bawt = dma_read_ctrl_rsci_biwt | dma_read_ctrl_rsci_bcwt;
  assign dma_read_ctrl_rsci_irdy_mxwt = MUX_s_1_2_2(dma_read_ctrl_rsci_irdy, dma_read_ctrl_rsci_irdy_bfwt,
      dma_read_ctrl_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_rsci_bcwt <= ~((~(dma_read_ctrl_rsci_bcwt | dma_read_ctrl_rsci_biwt))
          | dma_read_ctrl_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_irdy_bfwt <= 1'b0;
    end
    else if ( dma_read_ctrl_rsci_biwt ) begin
      dma_read_ctrl_rsci_irdy_bfwt <= dma_read_ctrl_rsci_irdy;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
    (
  core_wen, core_wten, dma_read_ctrl_rsci_oswt_unreg, dma_read_ctrl_rsci_iswt0, dma_read_ctrl_rsci_biwt,
      dma_read_ctrl_rsci_bdwt
);
  input core_wen;
  input core_wten;
  input dma_read_ctrl_rsci_oswt_unreg;
  input dma_read_ctrl_rsci_iswt0;
  output dma_read_ctrl_rsci_biwt;
  output dma_read_ctrl_rsci_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_rsci_bdwt = dma_read_ctrl_rsci_oswt_unreg & core_wen;
  assign dma_read_ctrl_rsci_biwt = (~ core_wten) & dma_read_ctrl_rsci_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp
    (
  clk, rst, plm_filters_rsci_bawt, plm_filters_rsci_biwt, plm_filters_rsci_bdwt
);
  input clk;
  input rst;
  output plm_filters_rsci_bawt;
  input plm_filters_rsci_biwt;
  input plm_filters_rsci_bdwt;


  // Interconnect Declarations
  reg plm_filters_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsci_bawt = plm_filters_rsci_biwt | plm_filters_rsci_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_filters_rsci_bcwt <= ~((~(plm_filters_rsci_bcwt | plm_filters_rsci_biwt))
          | plm_filters_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_filters_rsci_oswt_unreg, plm_filters_rsci_iswt0, plm_filters_rsci_biwt,
      plm_filters_rsci_bdwt, plm_filters_rsci_we_d_core_sct_pff, plm_filters_rsci_iswt0_pff
);
  input core_wen;
  input core_wten;
  input plm_filters_rsci_oswt_unreg;
  input plm_filters_rsci_iswt0;
  output plm_filters_rsci_biwt;
  output plm_filters_rsci_bdwt;
  output plm_filters_rsci_we_d_core_sct_pff;
  input plm_filters_rsci_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsci_bdwt = plm_filters_rsci_oswt_unreg & core_wen;
  assign plm_filters_rsci_biwt = (~ core_wten) & plm_filters_rsci_iswt0;
  assign plm_filters_rsci_we_d_core_sct_pff = plm_filters_rsci_iswt0_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp
    (
  clk, rst, plm_inputs_rsci_bawt, plm_inputs_rsci_biwt, plm_inputs_rsci_bdwt
);
  input clk;
  input rst;
  output plm_inputs_rsci_bawt;
  input plm_inputs_rsci_biwt;
  input plm_inputs_rsci_bdwt;


  // Interconnect Declarations
  reg plm_inputs_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsci_bawt = plm_inputs_rsci_biwt | plm_inputs_rsci_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_inputs_rsci_bcwt <= ~((~(plm_inputs_rsci_bcwt | plm_inputs_rsci_biwt))
          | plm_inputs_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_inputs_rsci_oswt_unreg, plm_inputs_rsci_iswt0, plm_inputs_rsci_biwt,
      plm_inputs_rsci_bdwt, plm_inputs_rsci_we_d_core_sct_pff, plm_inputs_rsci_iswt0_pff
);
  input core_wen;
  input core_wten;
  input plm_inputs_rsci_oswt_unreg;
  input plm_inputs_rsci_iswt0;
  output plm_inputs_rsci_biwt;
  output plm_inputs_rsci_bdwt;
  output plm_inputs_rsci_we_d_core_sct_pff;
  input plm_inputs_rsci_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsci_bdwt = plm_inputs_rsci_oswt_unreg & core_wen;
  assign plm_inputs_rsci_biwt = (~ core_wten) & plm_inputs_rsci_iswt0;
  assign plm_inputs_rsci_we_d_core_sct_pff = plm_inputs_rsci_iswt0_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_dp (
  clk, rst, conf_info_rsci_oswt_unreg, conf_info_rsci_bawt, conf_info_rsci_wen_comp,
      conf_info_rsci_idat_mxwt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  wire [231:0] conf_info_rsci_idat_mxwt_pconst;
  reg [231:0] conf_info_rsci_idat_bfwt_231_0;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bawt = conf_info_rsci_biwt | conf_info_rsci_bcwt;
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt_unreg) | conf_info_rsci_bawt;
  assign conf_info_rsci_idat_mxwt_pconst = MUX_v_232_2_2((conf_info_rsci_idat[231:0]),
      conf_info_rsci_idat_bfwt_231_0, conf_info_rsci_bcwt);
  assign conf_info_rsci_idat_mxwt = {(conf_info_rsci_idat_mxwt_pconst[231:224]) ,
      (conf_info_rsci_idat_mxwt_pconst[199:192]) , (conf_info_rsci_idat_mxwt_pconst[167:160])
      , (conf_info_rsci_idat_mxwt_pconst[135:128]) , (conf_info_rsci_idat_mxwt_pconst[103:96])
      , (conf_info_rsci_idat_mxwt_pconst[71:64]) , (conf_info_rsci_idat_mxwt_pconst[39:32])
      , (conf_info_rsci_idat_mxwt_pconst[7:0])};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt_231_0 <= conf_info_rsci_idat[231:0];
    end
  end

  function automatic [231:0] MUX_v_232_2_2;
    input [231:0] input_0;
    input [231:0] input_1;
    input [0:0] sel;
    reg [231:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_232_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_ctrl (
  core_wen, conf_info_rsci_oswt_unreg, conf_info_rsci_iswt0, conf_info_rsci_biwt,
      conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt_unreg & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_iswt0 & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_17_14_32_10368_10368_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_17_14_32_10368_10368_32_1_gen
    (
  we, d, wadr, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_16_32_50176_50176_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_16_32_50176_50176_32_1_gen
    (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [15:0] radr;
  output [31:0] q_d;
  input [15:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_15_14_32_10368_10368_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_15_14_32_10368_10368_32_1_gen
    (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output [31:0] q_d;
  input [13:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2d_cxx_catapult_compute_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2d_cxx_catapult_compute_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_staller (
  clk, rst, core_wen, core_wten, conf_info_rsci_wen_comp, done_rsci_wen_comp, plm_filters_rsc_req_obj_wen_comp,
      plm_inputs_rsc_req_obj_wen_comp, plm_outputs_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input conf_info_rsci_wen_comp;
  input done_rsci_wen_comp;
  input plm_filters_rsc_req_obj_wen_comp;
  input plm_inputs_rsc_req_obj_wen_comp;
  input plm_outputs_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & done_rsci_wen_comp & plm_filters_rsc_req_obj_wen_comp
      & plm_inputs_rsc_req_obj_wen_comp & plm_outputs_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp
    (
  clk, rst, plm_outputs_rsc_req_obj_oswt_unreg, plm_outputs_rsc_req_obj_bawt, plm_outputs_rsc_req_obj_wen_comp,
      plm_outputs_rsc_req_obj_biwt, plm_outputs_rsc_req_obj_bdwt, plm_outputs_rsc_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_outputs_rsc_req_obj_oswt_unreg;
  output plm_outputs_rsc_req_obj_bawt;
  output plm_outputs_rsc_req_obj_wen_comp;
  input plm_outputs_rsc_req_obj_biwt;
  input plm_outputs_rsc_req_obj_bdwt;
  output plm_outputs_rsc_req_obj_bcwt;
  reg plm_outputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_req_obj_bawt = plm_outputs_rsc_req_obj_biwt | plm_outputs_rsc_req_obj_bcwt;
  assign plm_outputs_rsc_req_obj_wen_comp = (~ plm_outputs_rsc_req_obj_oswt_unreg)
      | plm_outputs_rsc_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_outputs_rsc_req_obj_bcwt <= ~((~(plm_outputs_rsc_req_obj_bcwt | plm_outputs_rsc_req_obj_biwt))
          | plm_outputs_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl
    (
  core_wen, plm_outputs_rsc_req_obj_oswt_unreg, plm_outputs_rsc_req_obj_iswt0, plm_outputs_rsc_req_obj_vd,
      plm_outputs_rsc_req_obj_biwt, plm_outputs_rsc_req_obj_bdwt, plm_outputs_rsc_req_obj_bcwt
);
  input core_wen;
  input plm_outputs_rsc_req_obj_oswt_unreg;
  input plm_outputs_rsc_req_obj_iswt0;
  input plm_outputs_rsc_req_obj_vd;
  output plm_outputs_rsc_req_obj_biwt;
  output plm_outputs_rsc_req_obj_bdwt;
  input plm_outputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_req_obj_bdwt = plm_outputs_rsc_req_obj_oswt_unreg & core_wen;
  assign plm_outputs_rsc_req_obj_biwt = plm_outputs_rsc_req_obj_iswt0 & (~ plm_outputs_rsc_req_obj_bcwt)
      & plm_outputs_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp
    (
  clk, rst, plm_inputs_rsc_req_obj_oswt_unreg, plm_inputs_rsc_req_obj_bawt, plm_inputs_rsc_req_obj_wen_comp,
      plm_inputs_rsc_req_obj_biwt, plm_inputs_rsc_req_obj_bdwt, plm_inputs_rsc_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_inputs_rsc_req_obj_oswt_unreg;
  output plm_inputs_rsc_req_obj_bawt;
  output plm_inputs_rsc_req_obj_wen_comp;
  input plm_inputs_rsc_req_obj_biwt;
  input plm_inputs_rsc_req_obj_bdwt;
  output plm_inputs_rsc_req_obj_bcwt;
  reg plm_inputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_req_obj_bawt = plm_inputs_rsc_req_obj_biwt | plm_inputs_rsc_req_obj_bcwt;
  assign plm_inputs_rsc_req_obj_wen_comp = (~ plm_inputs_rsc_req_obj_oswt_unreg)
      | plm_inputs_rsc_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_inputs_rsc_req_obj_bcwt <= ~((~(plm_inputs_rsc_req_obj_bcwt | plm_inputs_rsc_req_obj_biwt))
          | plm_inputs_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl
    (
  core_wen, plm_inputs_rsc_req_obj_oswt_unreg, plm_inputs_rsc_req_obj_iswt0, plm_inputs_rsc_req_obj_vd,
      plm_inputs_rsc_req_obj_biwt, plm_inputs_rsc_req_obj_bdwt, plm_inputs_rsc_req_obj_bcwt
);
  input core_wen;
  input plm_inputs_rsc_req_obj_oswt_unreg;
  input plm_inputs_rsc_req_obj_iswt0;
  input plm_inputs_rsc_req_obj_vd;
  output plm_inputs_rsc_req_obj_biwt;
  output plm_inputs_rsc_req_obj_bdwt;
  input plm_inputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_req_obj_bdwt = plm_inputs_rsc_req_obj_oswt_unreg & core_wen;
  assign plm_inputs_rsc_req_obj_biwt = plm_inputs_rsc_req_obj_iswt0 & (~ plm_inputs_rsc_req_obj_bcwt)
      & plm_inputs_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp
    (
  clk, rst, plm_filters_rsc_req_obj_oswt_unreg, plm_filters_rsc_req_obj_bawt, plm_filters_rsc_req_obj_wen_comp,
      plm_filters_rsc_req_obj_biwt, plm_filters_rsc_req_obj_bdwt, plm_filters_rsc_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_filters_rsc_req_obj_oswt_unreg;
  output plm_filters_rsc_req_obj_bawt;
  output plm_filters_rsc_req_obj_wen_comp;
  input plm_filters_rsc_req_obj_biwt;
  input plm_filters_rsc_req_obj_bdwt;
  output plm_filters_rsc_req_obj_bcwt;
  reg plm_filters_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_req_obj_bawt = plm_filters_rsc_req_obj_biwt | plm_filters_rsc_req_obj_bcwt;
  assign plm_filters_rsc_req_obj_wen_comp = (~ plm_filters_rsc_req_obj_oswt_unreg)
      | plm_filters_rsc_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_filters_rsc_req_obj_bcwt <= ~((~(plm_filters_rsc_req_obj_bcwt | plm_filters_rsc_req_obj_biwt))
          | plm_filters_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl
    (
  core_wen, plm_filters_rsc_req_obj_oswt_unreg, plm_filters_rsc_req_obj_iswt0, plm_filters_rsc_req_obj_vd,
      plm_filters_rsc_req_obj_biwt, plm_filters_rsc_req_obj_bdwt, plm_filters_rsc_req_obj_bcwt
);
  input core_wen;
  input plm_filters_rsc_req_obj_oswt_unreg;
  input plm_filters_rsc_req_obj_iswt0;
  input plm_filters_rsc_req_obj_vd;
  output plm_filters_rsc_req_obj_biwt;
  output plm_filters_rsc_req_obj_bdwt;
  input plm_filters_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_req_obj_bdwt = plm_filters_rsc_req_obj_oswt_unreg & core_wen;
  assign plm_filters_rsc_req_obj_biwt = plm_filters_rsc_req_obj_iswt0 & (~ plm_filters_rsc_req_obj_bcwt)
      & plm_filters_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp
    (
  clk, rst, plm_filters_rsc_rls_obj_bawt, plm_filters_rsc_rls_obj_biwt, plm_filters_rsc_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_filters_rsc_rls_obj_bawt;
  input plm_filters_rsc_rls_obj_biwt;
  input plm_filters_rsc_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_filters_rsc_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_rls_obj_bawt = plm_filters_rsc_rls_obj_biwt | plm_filters_rsc_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsc_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_filters_rsc_rls_obj_bcwt <= ~((~(plm_filters_rsc_rls_obj_bcwt | plm_filters_rsc_rls_obj_biwt))
          | plm_filters_rsc_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl
    (
  core_wen, core_wten, plm_filters_rsc_rls_obj_oswt_unreg, plm_filters_rsc_rls_obj_iswt0,
      plm_filters_rsc_rls_obj_biwt, plm_filters_rsc_rls_obj_bdwt
);
  input core_wen;
  input core_wten;
  input plm_filters_rsc_rls_obj_oswt_unreg;
  input plm_filters_rsc_rls_obj_iswt0;
  output plm_filters_rsc_rls_obj_biwt;
  output plm_filters_rsc_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsc_rls_obj_bdwt = plm_filters_rsc_rls_obj_oswt_unreg & core_wen;
  assign plm_filters_rsc_rls_obj_biwt = (~ core_wten) & plm_filters_rsc_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp
    (
  clk, rst, plm_inputs_rsc_rls_obj_bawt, plm_inputs_rsc_rls_obj_biwt, plm_inputs_rsc_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_inputs_rsc_rls_obj_bawt;
  input plm_inputs_rsc_rls_obj_biwt;
  input plm_inputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_inputs_rsc_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_rls_obj_bawt = plm_inputs_rsc_rls_obj_biwt | plm_inputs_rsc_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsc_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_inputs_rsc_rls_obj_bcwt <= ~((~(plm_inputs_rsc_rls_obj_bcwt | plm_inputs_rsc_rls_obj_biwt))
          | plm_inputs_rsc_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl
    (
  core_wen, core_wten, plm_inputs_rsc_rls_obj_oswt_unreg, plm_inputs_rsc_rls_obj_iswt0,
      plm_inputs_rsc_rls_obj_biwt, plm_inputs_rsc_rls_obj_bdwt
);
  input core_wen;
  input core_wten;
  input plm_inputs_rsc_rls_obj_oswt_unreg;
  input plm_inputs_rsc_rls_obj_iswt0;
  output plm_inputs_rsc_rls_obj_biwt;
  output plm_inputs_rsc_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsc_rls_obj_bdwt = plm_inputs_rsc_rls_obj_oswt_unreg & core_wen;
  assign plm_inputs_rsc_rls_obj_biwt = (~ core_wten) & plm_inputs_rsc_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp
    (
  clk, rst, plm_outputs_rsc_rls_obj_bawt, plm_outputs_rsc_rls_obj_biwt, plm_outputs_rsc_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_outputs_rsc_rls_obj_bawt;
  input plm_outputs_rsc_rls_obj_biwt;
  input plm_outputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_outputs_rsc_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_rls_obj_bawt = plm_outputs_rsc_rls_obj_biwt | plm_outputs_rsc_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsc_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_outputs_rsc_rls_obj_bcwt <= ~((~(plm_outputs_rsc_rls_obj_bcwt | plm_outputs_rsc_rls_obj_biwt))
          | plm_outputs_rsc_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl
    (
  core_wen, core_wten, plm_outputs_rsc_rls_obj_oswt_unreg, plm_outputs_rsc_rls_obj_iswt0,
      plm_outputs_rsc_rls_obj_biwt, plm_outputs_rsc_rls_obj_bdwt
);
  input core_wen;
  input core_wten;
  input plm_outputs_rsc_rls_obj_oswt_unreg;
  input plm_outputs_rsc_rls_obj_iswt0;
  output plm_outputs_rsc_rls_obj_biwt;
  output plm_outputs_rsc_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_rls_obj_bdwt = plm_outputs_rsc_rls_obj_oswt_unreg & core_wen;
  assign plm_outputs_rsc_rls_obj_biwt = (~ core_wten) & plm_outputs_rsc_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt_unreg, done_rsci_bawt, done_rsci_wen_comp, done_rsci_biwt,
      done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bawt = done_rsci_biwt | done_rsci_bcwt;
  assign done_rsci_wen_comp = (~ done_rsci_oswt_unreg) | done_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt_unreg, done_rsci_iswt0, done_rsci_biwt, done_rsci_bdwt,
      done_rsci_bcwt, done_rsci_ivld_core_sct, done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt_unreg;
  input done_rsci_iswt0;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt_unreg & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_iswt0 & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp
    (
  clk, rst, plm_outputs_rsci_bawt, plm_outputs_rsci_biwt, plm_outputs_rsci_bdwt
);
  input clk;
  input rst;
  output plm_outputs_rsci_bawt;
  input plm_outputs_rsci_biwt;
  input plm_outputs_rsci_bdwt;


  // Interconnect Declarations
  reg plm_outputs_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsci_bawt = plm_outputs_rsci_biwt | plm_outputs_rsci_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_outputs_rsci_bcwt <= ~((~(plm_outputs_rsci_bcwt | plm_outputs_rsci_biwt))
          | plm_outputs_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_outputs_rsci_oswt_unreg, plm_outputs_rsci_iswt0, plm_outputs_rsci_biwt,
      plm_outputs_rsci_bdwt, plm_outputs_rsci_we_d_core_sct_pff, plm_outputs_rsci_iswt0_pff
);
  input core_wen;
  input core_wten;
  input plm_outputs_rsci_oswt_unreg;
  input plm_outputs_rsci_iswt0;
  output plm_outputs_rsci_biwt;
  output plm_outputs_rsci_bdwt;
  output plm_outputs_rsci_we_d_core_sct_pff;
  input plm_outputs_rsci_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsci_bdwt = plm_outputs_rsci_oswt_unreg & core_wen;
  assign plm_outputs_rsci_biwt = (~ core_wten) & plm_outputs_rsci_iswt0;
  assign plm_outputs_rsci_we_d_core_sct_pff = plm_outputs_rsci_iswt0_pff & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp
    (
  clk, rst, plm_filters_rsci_q_d, plm_filters_rsci_bawt, plm_filters_rsci_q_d_mxwt,
      plm_filters_rsci_biwt, plm_filters_rsci_bdwt
);
  input clk;
  input rst;
  input [31:0] plm_filters_rsci_q_d;
  output plm_filters_rsci_bawt;
  output [31:0] plm_filters_rsci_q_d_mxwt;
  input plm_filters_rsci_biwt;
  input plm_filters_rsci_bdwt;


  // Interconnect Declarations
  reg plm_filters_rsci_bcwt;
  reg [31:0] plm_filters_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsci_bawt = plm_filters_rsci_biwt | plm_filters_rsci_bcwt;
  assign plm_filters_rsci_q_d_mxwt = MUX_v_32_2_2(plm_filters_rsci_q_d, plm_filters_rsci_q_d_bfwt,
      plm_filters_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_filters_rsci_bcwt <= ~((~(plm_filters_rsci_bcwt | plm_filters_rsci_biwt))
          | plm_filters_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsci_q_d_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( plm_filters_rsci_biwt ) begin
      plm_filters_rsci_q_d_bfwt <= plm_filters_rsci_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_filters_rsci_oswt_unreg, plm_filters_rsci_iswt0, plm_filters_rsci_biwt,
      plm_filters_rsci_bdwt, plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct,
      plm_filters_rsci_iswt0_pff
);
  input core_wen;
  input core_wten;
  input plm_filters_rsci_oswt_unreg;
  input plm_filters_rsci_iswt0;
  output plm_filters_rsci_biwt;
  output plm_filters_rsci_bdwt;
  output plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  input plm_filters_rsci_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_filters_rsci_bdwt = plm_filters_rsci_oswt_unreg & core_wen;
  assign plm_filters_rsci_biwt = (~ core_wten) & plm_filters_rsci_iswt0;
  assign plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct = plm_filters_rsci_iswt0_pff
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp
    (
  clk, rst, plm_inputs_rsci_q_d, plm_inputs_rsci_bawt, plm_inputs_rsci_q_d_mxwt,
      plm_inputs_rsci_biwt, plm_inputs_rsci_bdwt
);
  input clk;
  input rst;
  input [31:0] plm_inputs_rsci_q_d;
  output plm_inputs_rsci_bawt;
  output [31:0] plm_inputs_rsci_q_d_mxwt;
  input plm_inputs_rsci_biwt;
  input plm_inputs_rsci_bdwt;


  // Interconnect Declarations
  reg plm_inputs_rsci_bcwt;
  reg [31:0] plm_inputs_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsci_bawt = plm_inputs_rsci_biwt | plm_inputs_rsci_bcwt;
  assign plm_inputs_rsci_q_d_mxwt = MUX_v_32_2_2(plm_inputs_rsci_q_d, plm_inputs_rsci_q_d_bfwt,
      plm_inputs_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_inputs_rsci_bcwt <= ~((~(plm_inputs_rsci_bcwt | plm_inputs_rsci_biwt))
          | plm_inputs_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsci_q_d_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( plm_inputs_rsci_biwt ) begin
      plm_inputs_rsci_q_d_bfwt <= plm_inputs_rsci_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_inputs_rsci_oswt_unreg, plm_inputs_rsci_iswt0, plm_inputs_rsci_biwt,
      plm_inputs_rsci_bdwt, plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct,
      plm_inputs_rsci_iswt0_pff
);
  input core_wen;
  input core_wten;
  input plm_inputs_rsci_oswt_unreg;
  input plm_inputs_rsci_iswt0;
  output plm_inputs_rsci_biwt;
  output plm_inputs_rsci_bdwt;
  output plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  input plm_inputs_rsci_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_inputs_rsci_bdwt = plm_inputs_rsci_oswt_unreg & core_wen;
  assign plm_inputs_rsci_biwt = (~ core_wten) & plm_inputs_rsci_iswt0;
  assign plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct = plm_inputs_rsci_iswt0_pff
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_dp
    (
  clk, rst, conf_info_rsci_oswt_unreg, conf_info_rsci_bawt, conf_info_rsci_wen_comp,
      conf_info_rsci_idat_mxwt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  wire [231:0] conf_info_rsci_idat_mxwt_pconst;
  reg [231:0] conf_info_rsci_idat_bfwt_231_0;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bawt = conf_info_rsci_biwt | conf_info_rsci_bcwt;
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt_unreg) | conf_info_rsci_bawt;
  assign conf_info_rsci_idat_mxwt_pconst = MUX_v_232_2_2((conf_info_rsci_idat[231:0]),
      conf_info_rsci_idat_bfwt_231_0, conf_info_rsci_bcwt);
  assign conf_info_rsci_idat_mxwt = {(conf_info_rsci_idat_mxwt_pconst[231:224]) ,
      (conf_info_rsci_idat_mxwt_pconst[199:192]) , (conf_info_rsci_idat_mxwt_pconst[167:160])
      , (conf_info_rsci_idat_mxwt_pconst[135:128]) , (conf_info_rsci_idat_mxwt_pconst[103:96])
      , (conf_info_rsci_idat_mxwt_pconst[71:64]) , (conf_info_rsci_idat_mxwt_pconst[39:32])
      , (conf_info_rsci_idat_mxwt_pconst[7:0])};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt_231_0 <= conf_info_rsci_idat[231:0];
    end
  end

  function automatic [231:0] MUX_v_232_2_2;
    input [231:0] input_0;
    input [231:0] input_1;
    input [0:0] sel;
    reg [231:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_232_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt_unreg, conf_info_rsci_iswt0, conf_info_rsci_biwt,
      conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt_unreg & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_iswt0 & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_24_14_32_10368_10368_32_1_gen
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_24_14_32_10368_10368_32_1_gen
    (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output [31:0] q_d;
  input [13:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for esp_acc_conv2d_cxx_catapult_store_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_conv2d_cxx_catapult_store_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_staller
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_staller (
  clk, rst, core_wen, core_wten, conf_info_rsci_wen_comp, dma_write_ctrl_rsci_wen_comp,
      dma_write_chnl_rsci_wen_comp, done_rsci_wen_comp, plm_outputs_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  input conf_info_rsci_wen_comp;
  input dma_write_ctrl_rsci_wen_comp;
  input dma_write_chnl_rsci_wen_comp;
  input done_rsci_wen_comp;
  input plm_outputs_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = conf_info_rsci_wen_comp & dma_write_ctrl_rsci_wen_comp & dma_write_chnl_rsci_wen_comp
      & done_rsci_wen_comp & plm_outputs_rsc_req_obj_wen_comp;
  assign core_wten = core_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp
    (
  clk, rst, plm_outputs_rsc_req_obj_oswt_unreg, plm_outputs_rsc_req_obj_bawt, plm_outputs_rsc_req_obj_wen_comp,
      plm_outputs_rsc_req_obj_biwt, plm_outputs_rsc_req_obj_bdwt, plm_outputs_rsc_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_outputs_rsc_req_obj_oswt_unreg;
  output plm_outputs_rsc_req_obj_bawt;
  output plm_outputs_rsc_req_obj_wen_comp;
  input plm_outputs_rsc_req_obj_biwt;
  input plm_outputs_rsc_req_obj_bdwt;
  output plm_outputs_rsc_req_obj_bcwt;
  reg plm_outputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_req_obj_bawt = plm_outputs_rsc_req_obj_biwt | plm_outputs_rsc_req_obj_bcwt;
  assign plm_outputs_rsc_req_obj_wen_comp = (~ plm_outputs_rsc_req_obj_oswt_unreg)
      | plm_outputs_rsc_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_outputs_rsc_req_obj_bcwt <= ~((~(plm_outputs_rsc_req_obj_bcwt | plm_outputs_rsc_req_obj_biwt))
          | plm_outputs_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl
    (
  core_wen, plm_outputs_rsc_req_obj_oswt_unreg, plm_outputs_rsc_req_obj_iswt0, plm_outputs_rsc_req_obj_vd,
      plm_outputs_rsc_req_obj_biwt, plm_outputs_rsc_req_obj_bdwt, plm_outputs_rsc_req_obj_bcwt
);
  input core_wen;
  input plm_outputs_rsc_req_obj_oswt_unreg;
  input plm_outputs_rsc_req_obj_iswt0;
  input plm_outputs_rsc_req_obj_vd;
  output plm_outputs_rsc_req_obj_biwt;
  output plm_outputs_rsc_req_obj_bdwt;
  input plm_outputs_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_req_obj_bdwt = plm_outputs_rsc_req_obj_oswt_unreg & core_wen;
  assign plm_outputs_rsc_req_obj_biwt = plm_outputs_rsc_req_obj_iswt0 & (~ plm_outputs_rsc_req_obj_bcwt)
      & plm_outputs_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp
    (
  clk, rst, plm_outputs_rsc_rls_obj_bawt, plm_outputs_rsc_rls_obj_biwt, plm_outputs_rsc_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_outputs_rsc_rls_obj_bawt;
  input plm_outputs_rsc_rls_obj_biwt;
  input plm_outputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_outputs_rsc_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_rls_obj_bawt = plm_outputs_rsc_rls_obj_biwt | plm_outputs_rsc_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsc_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_outputs_rsc_rls_obj_bcwt <= ~((~(plm_outputs_rsc_rls_obj_bcwt | plm_outputs_rsc_rls_obj_biwt))
          | plm_outputs_rsc_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl
    (
  core_wen, core_wten, plm_outputs_rsc_rls_obj_oswt_unreg, plm_outputs_rsc_rls_obj_iswt0,
      plm_outputs_rsc_rls_obj_biwt, plm_outputs_rsc_rls_obj_bdwt
);
  input core_wen;
  input core_wten;
  input plm_outputs_rsc_rls_obj_oswt_unreg;
  input plm_outputs_rsc_rls_obj_iswt0;
  output plm_outputs_rsc_rls_obj_biwt;
  output plm_outputs_rsc_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsc_rls_obj_bdwt = plm_outputs_rsc_rls_obj_oswt_unreg & core_wen;
  assign plm_outputs_rsc_rls_obj_biwt = (~ core_wten) & plm_outputs_rsc_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_done_rsci_done_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_done_rsci_done_wait_dp (
  clk, rst, done_rsci_oswt_unreg, done_rsci_bawt, done_rsci_wen_comp, done_rsci_biwt,
      done_rsci_bdwt, done_rsci_bcwt
);
  input clk;
  input rst;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  output done_rsci_wen_comp;
  input done_rsci_biwt;
  input done_rsci_bdwt;
  output done_rsci_bcwt;
  reg done_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bawt = done_rsci_biwt | done_rsci_bcwt;
  assign done_rsci_wen_comp = (~ done_rsci_oswt_unreg) | done_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done_rsci_bcwt <= 1'b0;
    end
    else begin
      done_rsci_bcwt <= ~((~(done_rsci_bcwt | done_rsci_biwt)) | done_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_done_rsci_done_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_done_rsci_done_wait_ctrl (
  core_wen, done_rsci_oswt_unreg, done_rsci_iswt0, done_rsci_biwt, done_rsci_bdwt,
      done_rsci_bcwt, done_rsci_ivld_core_sct, done_rsci_irdy
);
  input core_wen;
  input done_rsci_oswt_unreg;
  input done_rsci_iswt0;
  output done_rsci_biwt;
  output done_rsci_bdwt;
  input done_rsci_bcwt;
  output done_rsci_ivld_core_sct;
  input done_rsci_irdy;


  // Interconnect Declarations
  wire done_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign done_rsci_bdwt = done_rsci_oswt_unreg & core_wen;
  assign done_rsci_biwt = done_rsci_ogwt & done_rsci_irdy;
  assign done_rsci_ogwt = done_rsci_iswt0 & (~ done_rsci_bcwt);
  assign done_rsci_ivld_core_sct = done_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
    (
  clk, rst, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_bawt, dma_write_chnl_rsci_wen_comp,
      dma_write_chnl_rsci_biwt, dma_write_chnl_rsci_bdwt, dma_write_chnl_rsci_bcwt
);
  input clk;
  input rst;
  input dma_write_chnl_rsci_oswt_unreg;
  output dma_write_chnl_rsci_bawt;
  output dma_write_chnl_rsci_wen_comp;
  input dma_write_chnl_rsci_biwt;
  input dma_write_chnl_rsci_bdwt;
  output dma_write_chnl_rsci_bcwt;
  reg dma_write_chnl_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_rsci_bawt = dma_write_chnl_rsci_biwt | dma_write_chnl_rsci_bcwt;
  assign dma_write_chnl_rsci_wen_comp = (~ dma_write_chnl_rsci_oswt_unreg) | dma_write_chnl_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_write_chnl_rsci_bcwt <= ~((~(dma_write_chnl_rsci_bcwt | dma_write_chnl_rsci_biwt))
          | dma_write_chnl_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
    (
  core_wen, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_iswt0, dma_write_chnl_rsci_irdy,
      dma_write_chnl_rsci_biwt, dma_write_chnl_rsci_bdwt, dma_write_chnl_rsci_bcwt,
      dma_write_chnl_rsci_ivld_core_sct
);
  input core_wen;
  input dma_write_chnl_rsci_oswt_unreg;
  input dma_write_chnl_rsci_iswt0;
  input dma_write_chnl_rsci_irdy;
  output dma_write_chnl_rsci_biwt;
  output dma_write_chnl_rsci_bdwt;
  input dma_write_chnl_rsci_bcwt;
  output dma_write_chnl_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire dma_write_chnl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_rsci_bdwt = dma_write_chnl_rsci_oswt_unreg & core_wen;
  assign dma_write_chnl_rsci_biwt = dma_write_chnl_rsci_ogwt & dma_write_chnl_rsci_irdy;
  assign dma_write_chnl_rsci_ogwt = dma_write_chnl_rsci_iswt0 & (~ dma_write_chnl_rsci_bcwt);
  assign dma_write_chnl_rsci_ivld_core_sct = dma_write_chnl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
    (
  clk, rst, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_bawt, dma_write_ctrl_rsci_wen_comp,
      dma_write_ctrl_rsci_biwt, dma_write_ctrl_rsci_bdwt, dma_write_ctrl_rsci_bcwt
);
  input clk;
  input rst;
  input dma_write_ctrl_rsci_oswt_unreg;
  output dma_write_ctrl_rsci_bawt;
  output dma_write_ctrl_rsci_wen_comp;
  input dma_write_ctrl_rsci_biwt;
  input dma_write_ctrl_rsci_bdwt;
  output dma_write_ctrl_rsci_bcwt;
  reg dma_write_ctrl_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_rsci_bawt = dma_write_ctrl_rsci_biwt | dma_write_ctrl_rsci_bcwt;
  assign dma_write_ctrl_rsci_wen_comp = (~ dma_write_ctrl_rsci_oswt_unreg) | dma_write_ctrl_rsci_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_rsci_bcwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_rsci_bcwt <= ~((~(dma_write_ctrl_rsci_bcwt | dma_write_ctrl_rsci_biwt))
          | dma_write_ctrl_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
    (
  core_wen, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_iswt0, dma_write_ctrl_rsci_irdy,
      dma_write_ctrl_rsci_biwt, dma_write_ctrl_rsci_bdwt, dma_write_ctrl_rsci_bcwt,
      dma_write_ctrl_rsci_ivld_core_sct
);
  input core_wen;
  input dma_write_ctrl_rsci_oswt_unreg;
  input dma_write_ctrl_rsci_iswt0;
  input dma_write_ctrl_rsci_irdy;
  output dma_write_ctrl_rsci_biwt;
  output dma_write_ctrl_rsci_bdwt;
  input dma_write_ctrl_rsci_bcwt;
  output dma_write_ctrl_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire dma_write_ctrl_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_rsci_bdwt = dma_write_ctrl_rsci_oswt_unreg & core_wen;
  assign dma_write_ctrl_rsci_biwt = dma_write_ctrl_rsci_ogwt & dma_write_ctrl_rsci_irdy;
  assign dma_write_ctrl_rsci_ogwt = dma_write_ctrl_rsci_iswt0 & (~ dma_write_ctrl_rsci_bcwt);
  assign dma_write_ctrl_rsci_ivld_core_sct = dma_write_ctrl_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp
    (
  clk, rst, plm_outputs_rsci_q_d, plm_outputs_rsci_bawt, plm_outputs_rsci_q_d_mxwt,
      plm_outputs_rsci_biwt, plm_outputs_rsci_bdwt
);
  input clk;
  input rst;
  input [31:0] plm_outputs_rsci_q_d;
  output plm_outputs_rsci_bawt;
  output [31:0] plm_outputs_rsci_q_d_mxwt;
  input plm_outputs_rsci_biwt;
  input plm_outputs_rsci_bdwt;


  // Interconnect Declarations
  reg plm_outputs_rsci_bcwt;
  reg [31:0] plm_outputs_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsci_bawt = plm_outputs_rsci_biwt | plm_outputs_rsci_bcwt;
  assign plm_outputs_rsci_q_d_mxwt = MUX_v_32_2_2(plm_outputs_rsci_q_d, plm_outputs_rsci_q_d_bfwt,
      plm_outputs_rsci_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsci_bcwt <= 1'b0;
    end
    else begin
      plm_outputs_rsci_bcwt <= ~((~(plm_outputs_rsci_bcwt | plm_outputs_rsci_biwt))
          | plm_outputs_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsci_q_d_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( plm_outputs_rsci_biwt ) begin
      plm_outputs_rsci_q_d_bfwt <= plm_outputs_rsci_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl
    (
  core_wen, core_wten, plm_outputs_rsci_oswt_unreg, plm_outputs_rsci_iswt0, plm_outputs_rsci_biwt,
      plm_outputs_rsci_bdwt, plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct,
      plm_outputs_rsci_iswt0_pff
);
  input core_wen;
  input core_wten;
  input plm_outputs_rsci_oswt_unreg;
  input plm_outputs_rsci_iswt0;
  output plm_outputs_rsci_biwt;
  output plm_outputs_rsci_bdwt;
  output plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
  input plm_outputs_rsci_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_outputs_rsci_bdwt = plm_outputs_rsci_oswt_unreg & core_wen;
  assign plm_outputs_rsci_biwt = (~ core_wten) & plm_outputs_rsci_iswt0;
  assign plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct = plm_outputs_rsci_iswt0_pff
      & core_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_dp
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_dp (
  clk, rst, conf_info_rsci_oswt_unreg, conf_info_rsci_bawt, conf_info_rsci_wen_comp,
      conf_info_rsci_idat_mxwt, conf_info_rsci_biwt, conf_info_rsci_bdwt, conf_info_rsci_bcwt,
      conf_info_rsci_idat
);
  input clk;
  input rst;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;
  input conf_info_rsci_biwt;
  input conf_info_rsci_bdwt;
  output conf_info_rsci_bcwt;
  reg conf_info_rsci_bcwt;
  input [255:0] conf_info_rsci_idat;


  // Interconnect Declarations
  wire [231:0] conf_info_rsci_idat_mxwt_pconst;
  reg [231:0] conf_info_rsci_idat_bfwt_231_0;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bawt = conf_info_rsci_biwt | conf_info_rsci_bcwt;
  assign conf_info_rsci_wen_comp = (~ conf_info_rsci_oswt_unreg) | conf_info_rsci_bawt;
  assign conf_info_rsci_idat_mxwt_pconst = MUX_v_232_2_2((conf_info_rsci_idat[231:0]),
      conf_info_rsci_idat_bfwt_231_0, conf_info_rsci_bcwt);
  assign conf_info_rsci_idat_mxwt = {(conf_info_rsci_idat_mxwt_pconst[231:224]) ,
      (conf_info_rsci_idat_mxwt_pconst[199:192]) , (conf_info_rsci_idat_mxwt_pconst[167:160])
      , (conf_info_rsci_idat_mxwt_pconst[135:128]) , (conf_info_rsci_idat_mxwt_pconst[103:96])
      , (conf_info_rsci_idat_mxwt_pconst[71:64]) , (conf_info_rsci_idat_mxwt_pconst[39:32])
      , (conf_info_rsci_idat_mxwt_pconst[7:0])};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_bcwt <= 1'b0;
    end
    else begin
      conf_info_rsci_bcwt <= ~((~(conf_info_rsci_bcwt | conf_info_rsci_biwt)) | conf_info_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      conf_info_rsci_idat_bfwt_231_0 <= 232'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( conf_info_rsci_biwt ) begin
      conf_info_rsci_idat_bfwt_231_0 <= conf_info_rsci_idat[231:0];
    end
  end

  function automatic [231:0] MUX_v_232_2_2;
    input [231:0] input_0;
    input [231:0] input_1;
    input [0:0] sel;
    reg [231:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_232_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_ctrl
    (
  core_wen, conf_info_rsci_oswt_unreg, conf_info_rsci_iswt0, conf_info_rsci_biwt,
      conf_info_rsci_bdwt, conf_info_rsci_bcwt, conf_info_rsci_irdy_core_sct, conf_info_rsci_ivld
);
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_biwt;
  output conf_info_rsci_bdwt;
  input conf_info_rsci_bcwt;
  output conf_info_rsci_irdy_core_sct;
  input conf_info_rsci_ivld;


  // Interconnect Declarations
  wire conf_info_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign conf_info_rsci_bdwt = conf_info_rsci_oswt_unreg & core_wen;
  assign conf_info_rsci_biwt = conf_info_rsci_ogwt & conf_info_rsci_ivld;
  assign conf_info_rsci_ogwt = conf_info_rsci_iswt0 & (~ conf_info_rsci_bcwt);
  assign conf_info_rsci_irdy_core_sct = conf_info_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi
    (
  clk, rst, store_done_cns_rdy, store_done_cns_vld, core_wen, store_done_cnsi_oswt_unreg,
      store_done_cnsi_bawt, store_done_cnsi_iswt0, store_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output store_done_cns_rdy;
  input store_done_cns_vld;
  input core_wen;
  input store_done_cnsi_oswt_unreg;
  output store_done_cnsi_bawt;
  input store_done_cnsi_iswt0;
  output store_done_cnsi_wen_comp;


  // Interconnect Declarations
  wire store_done_cnsi_ivld;
  wire store_done_cnsi_biwt;
  wire store_done_cnsi_bdwt;
  wire store_done_cnsi_bcwt;
  wire store_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd49)) store_done_cnsi
      (
      .vld(store_done_cns_vld),
      .rdy(store_done_cns_rdy),
      .ivld(store_done_cnsi_ivld),
      .irdy(store_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl
      conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_ctrl_inst (
      .core_wen(core_wen),
      .store_done_cnsi_oswt_unreg(store_done_cnsi_oswt_unreg),
      .store_done_cnsi_iswt0(store_done_cnsi_iswt0),
      .store_done_cnsi_ivld(store_done_cnsi_ivld),
      .store_done_cnsi_biwt(store_done_cnsi_biwt),
      .store_done_cnsi_bdwt(store_done_cnsi_bdwt),
      .store_done_cnsi_bcwt(store_done_cnsi_bcwt),
      .store_done_cnsi_irdy_core_sct(store_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp
      conv2d_cxx_catapult_core_core_store_done_cnsi_store_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .store_done_cnsi_oswt_unreg(store_done_cnsi_oswt_unreg),
      .store_done_cnsi_bawt(store_done_cnsi_bawt),
      .store_done_cnsi_wen_comp(store_done_cnsi_wen_comp),
      .store_done_cnsi_biwt(store_done_cnsi_biwt),
      .store_done_cnsi_bdwt(store_done_cnsi_bdwt),
      .store_done_cnsi_bcwt(store_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi
    (
  clk, rst, compute_done_cns_rdy, compute_done_cns_vld, core_wen, compute_done_cnsi_oswt_unreg,
      compute_done_cnsi_bawt, compute_done_cnsi_iswt0, compute_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output compute_done_cns_rdy;
  input compute_done_cns_vld;
  input core_wen;
  input compute_done_cnsi_oswt_unreg;
  output compute_done_cnsi_bawt;
  input compute_done_cnsi_iswt0;
  output compute_done_cnsi_wen_comp;


  // Interconnect Declarations
  wire compute_done_cnsi_ivld;
  wire compute_done_cnsi_biwt;
  wire compute_done_cnsi_bdwt;
  wire compute_done_cnsi_bcwt;
  wire compute_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd48)) compute_done_cnsi
      (
      .vld(compute_done_cns_vld),
      .rdy(compute_done_cns_rdy),
      .ivld(compute_done_cnsi_ivld),
      .irdy(compute_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl
      conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .compute_done_cnsi_oswt_unreg(compute_done_cnsi_oswt_unreg),
      .compute_done_cnsi_iswt0(compute_done_cnsi_iswt0),
      .compute_done_cnsi_ivld(compute_done_cnsi_ivld),
      .compute_done_cnsi_biwt(compute_done_cnsi_biwt),
      .compute_done_cnsi_bdwt(compute_done_cnsi_bdwt),
      .compute_done_cnsi_bcwt(compute_done_cnsi_bcwt),
      .compute_done_cnsi_irdy_core_sct(compute_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp
      conv2d_cxx_catapult_core_core_compute_done_cnsi_compute_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .compute_done_cnsi_oswt_unreg(compute_done_cnsi_oswt_unreg),
      .compute_done_cnsi_bawt(compute_done_cnsi_bawt),
      .compute_done_cnsi_wen_comp(compute_done_cnsi_wen_comp),
      .compute_done_cnsi_biwt(compute_done_cnsi_biwt),
      .compute_done_cnsi_bdwt(compute_done_cnsi_bdwt),
      .compute_done_cnsi_bcwt(compute_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi (
  clk, rst, load_done_cns_rdy, load_done_cns_vld, core_wen, load_done_cnsi_oswt_unreg,
      load_done_cnsi_bawt, load_done_cnsi_iswt0, load_done_cnsi_wen_comp, load_done_cnsi_irdy_core_psct
);
  input clk;
  input rst;
  output load_done_cns_rdy;
  input load_done_cns_vld;
  input core_wen;
  input load_done_cnsi_oswt_unreg;
  output load_done_cnsi_bawt;
  input load_done_cnsi_iswt0;
  output load_done_cnsi_wen_comp;
  input load_done_cnsi_irdy_core_psct;


  // Interconnect Declarations
  wire load_done_cnsi_ivld;
  wire load_done_cnsi_biwt;
  wire load_done_cnsi_bdwt;
  wire load_done_cnsi_bcwt;
  wire load_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd47)) load_done_cnsi
      (
      .vld(load_done_cns_vld),
      .rdy(load_done_cns_rdy),
      .ivld(load_done_cnsi_ivld),
      .irdy(load_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl
      conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_ctrl_inst (
      .core_wen(core_wen),
      .load_done_cnsi_oswt_unreg(load_done_cnsi_oswt_unreg),
      .load_done_cnsi_iswt0(load_done_cnsi_iswt0),
      .load_done_cnsi_irdy_core_psct(load_done_cnsi_irdy_core_psct),
      .load_done_cnsi_ivld(load_done_cnsi_ivld),
      .load_done_cnsi_biwt(load_done_cnsi_biwt),
      .load_done_cnsi_bdwt(load_done_cnsi_bdwt),
      .load_done_cnsi_bcwt(load_done_cnsi_bcwt),
      .load_done_cnsi_irdy_core_sct(load_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp
      conv2d_cxx_catapult_core_core_load_done_cnsi_load_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .load_done_cnsi_oswt_unreg(load_done_cnsi_oswt_unreg),
      .load_done_cnsi_bawt(load_done_cnsi_bawt),
      .load_done_cnsi_wen_comp(load_done_cnsi_wen_comp),
      .load_done_cnsi_biwt(load_done_cnsi_biwt),
      .load_done_cnsi_bdwt(load_done_cnsi_bdwt),
      .load_done_cnsi_bcwt(load_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi
    (
  clk, rst, config_done_cns_rdy, config_done_cns_vld, core_wen, config_done_cnsi_oswt_unreg,
      config_done_cnsi_bawt, config_done_cnsi_iswt0, config_done_cnsi_wen_comp
);
  input clk;
  input rst;
  output config_done_cns_rdy;
  input config_done_cns_vld;
  input core_wen;
  input config_done_cnsi_oswt_unreg;
  output config_done_cnsi_bawt;
  input config_done_cnsi_iswt0;
  output config_done_cnsi_wen_comp;


  // Interconnect Declarations
  wire config_done_cnsi_ivld;
  wire config_done_cnsi_biwt;
  wire config_done_cnsi_bdwt;
  wire config_done_cnsi_bcwt;
  wire config_done_cnsi_irdy_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_in_wait_v1 #(.rscid(32'sd46)) config_done_cnsi
      (
      .vld(config_done_cns_vld),
      .rdy(config_done_cns_rdy),
      .ivld(config_done_cnsi_ivld),
      .irdy(config_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl
      conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_ctrl_inst (
      .core_wen(core_wen),
      .config_done_cnsi_oswt_unreg(config_done_cnsi_oswt_unreg),
      .config_done_cnsi_iswt0(config_done_cnsi_iswt0),
      .config_done_cnsi_ivld(config_done_cnsi_ivld),
      .config_done_cnsi_biwt(config_done_cnsi_biwt),
      .config_done_cnsi_bdwt(config_done_cnsi_bdwt),
      .config_done_cnsi_bcwt(config_done_cnsi_bcwt),
      .config_done_cnsi_irdy_core_sct(config_done_cnsi_irdy_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp
      conv2d_cxx_catapult_core_core_config_done_cnsi_config_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .config_done_cnsi_oswt_unreg(config_done_cnsi_oswt_unreg),
      .config_done_cnsi_bawt(config_done_cnsi_bawt),
      .config_done_cnsi_wen_comp(config_done_cnsi_wen_comp),
      .config_done_cnsi_biwt(config_done_cnsi_biwt),
      .config_done_cnsi_bdwt(config_done_cnsi_bdwt),
      .config_done_cnsi_bcwt(config_done_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci (
  clk, rst, acc_done_rsc_vld, core_wen, acc_done_rsci_oswt_unreg, acc_done_rsci_bawt,
      acc_done_rsci_iswt0, core_wten
);
  input clk;
  input rst;
  output acc_done_rsc_vld;
  input core_wen;
  input acc_done_rsci_oswt_unreg;
  output acc_done_rsci_bawt;
  input acc_done_rsci_iswt0;
  input core_wten;


  // Interconnect Declarations
  wire acc_done_rsci_biwt;
  wire acc_done_rsci_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_out_vld_v1 #(.rscid(32'sd45)) acc_done_rsci
      (
      .vld(acc_done_rsc_vld),
      .ivld(acc_done_rsci_biwt)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl
      conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_ctrl_inst (
      .core_wen(core_wen),
      .acc_done_rsci_oswt_unreg(acc_done_rsci_oswt_unreg),
      .acc_done_rsci_iswt0(acc_done_rsci_iswt0),
      .core_wten(core_wten),
      .acc_done_rsci_biwt(acc_done_rsci_biwt),
      .acc_done_rsci_bdwt(acc_done_rsci_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp
      conv2d_cxx_catapult_core_core_acc_done_rsci_acc_done_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .acc_done_rsci_bawt(acc_done_rsci_bawt),
      .acc_done_rsci_biwt(acc_done_rsci_biwt),
      .acc_done_rsci_bdwt(acc_done_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt_unreg, done_rsci_bawt,
      done_rsci_iswt0, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  input done_rsci_iswt0;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd5)) done_rsci (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_config_core_done_rsci_done_wait_ctrl config_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_iswt0(done_rsci_iswt0),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_config_core_done_rsci_done_wait_dp config_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci (
  clk, rst, plm_conf_store_rsc_dat, plm_conf_store_rsc_vld, plm_conf_store_rsc_rdy,
      core_wen, plm_conf_store_rsci_oswt_unreg, plm_conf_store_rsci_bawt, plm_conf_store_rsci_iswt0,
      plm_conf_store_rsci_wen_comp, plm_conf_store_rsci_idat
);
  input clk;
  input rst;
  output [255:0] plm_conf_store_rsc_dat;
  output plm_conf_store_rsc_vld;
  input plm_conf_store_rsc_rdy;
  input core_wen;
  input plm_conf_store_rsci_oswt_unreg;
  output plm_conf_store_rsci_bawt;
  input plm_conf_store_rsci_iswt0;
  output plm_conf_store_rsci_wen_comp;
  input [255:0] plm_conf_store_rsci_idat;


  // Interconnect Declarations
  wire plm_conf_store_rsci_irdy;
  wire plm_conf_store_rsci_biwt;
  wire plm_conf_store_rsci_bdwt;
  wire plm_conf_store_rsci_bcwt;
  wire plm_conf_store_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd256)) plm_conf_store_rsci (
      .irdy(plm_conf_store_rsci_irdy),
      .ivld(plm_conf_store_rsci_ivld_core_sct),
      .idat(plm_conf_store_rsci_idat),
      .rdy(plm_conf_store_rsc_rdy),
      .vld(plm_conf_store_rsc_vld),
      .dat(plm_conf_store_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl
      config_core_plm_conf_store_rsci_plm_conf_store_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_conf_store_rsci_oswt_unreg(plm_conf_store_rsci_oswt_unreg),
      .plm_conf_store_rsci_iswt0(plm_conf_store_rsci_iswt0),
      .plm_conf_store_rsci_irdy(plm_conf_store_rsci_irdy),
      .plm_conf_store_rsci_biwt(plm_conf_store_rsci_biwt),
      .plm_conf_store_rsci_bdwt(plm_conf_store_rsci_bdwt),
      .plm_conf_store_rsci_bcwt(plm_conf_store_rsci_bcwt),
      .plm_conf_store_rsci_ivld_core_sct(plm_conf_store_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci_plm_conf_store_wait_dp
      config_core_plm_conf_store_rsci_plm_conf_store_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_conf_store_rsci_oswt_unreg(plm_conf_store_rsci_oswt_unreg),
      .plm_conf_store_rsci_bawt(plm_conf_store_rsci_bawt),
      .plm_conf_store_rsci_wen_comp(plm_conf_store_rsci_wen_comp),
      .plm_conf_store_rsci_biwt(plm_conf_store_rsci_biwt),
      .plm_conf_store_rsci_bdwt(plm_conf_store_rsci_bdwt),
      .plm_conf_store_rsci_bcwt(plm_conf_store_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci (
  clk, rst, plm_conf_compute_rsc_dat, plm_conf_compute_rsc_vld, plm_conf_compute_rsc_rdy,
      core_wen, plm_conf_compute_rsci_oswt_unreg, plm_conf_compute_rsci_bawt, plm_conf_compute_rsci_iswt0,
      plm_conf_compute_rsci_wen_comp, plm_conf_compute_rsci_idat
);
  input clk;
  input rst;
  output [255:0] plm_conf_compute_rsc_dat;
  output plm_conf_compute_rsc_vld;
  input plm_conf_compute_rsc_rdy;
  input core_wen;
  input plm_conf_compute_rsci_oswt_unreg;
  output plm_conf_compute_rsci_bawt;
  input plm_conf_compute_rsci_iswt0;
  output plm_conf_compute_rsci_wen_comp;
  input [255:0] plm_conf_compute_rsci_idat;


  // Interconnect Declarations
  wire plm_conf_compute_rsci_irdy;
  wire plm_conf_compute_rsci_biwt;
  wire plm_conf_compute_rsci_bdwt;
  wire plm_conf_compute_rsci_bcwt;
  wire plm_conf_compute_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd256)) plm_conf_compute_rsci (
      .irdy(plm_conf_compute_rsci_irdy),
      .ivld(plm_conf_compute_rsci_ivld_core_sct),
      .idat(plm_conf_compute_rsci_idat),
      .rdy(plm_conf_compute_rsc_rdy),
      .vld(plm_conf_compute_rsc_vld),
      .dat(plm_conf_compute_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl
      config_core_plm_conf_compute_rsci_plm_conf_compute_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_conf_compute_rsci_oswt_unreg(plm_conf_compute_rsci_oswt_unreg),
      .plm_conf_compute_rsci_iswt0(plm_conf_compute_rsci_iswt0),
      .plm_conf_compute_rsci_irdy(plm_conf_compute_rsci_irdy),
      .plm_conf_compute_rsci_biwt(plm_conf_compute_rsci_biwt),
      .plm_conf_compute_rsci_bdwt(plm_conf_compute_rsci_bdwt),
      .plm_conf_compute_rsci_bcwt(plm_conf_compute_rsci_bcwt),
      .plm_conf_compute_rsci_ivld_core_sct(plm_conf_compute_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp
      config_core_plm_conf_compute_rsci_plm_conf_compute_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_conf_compute_rsci_oswt_unreg(plm_conf_compute_rsci_oswt_unreg),
      .plm_conf_compute_rsci_bawt(plm_conf_compute_rsci_bawt),
      .plm_conf_compute_rsci_wen_comp(plm_conf_compute_rsci_wen_comp),
      .plm_conf_compute_rsci_biwt(plm_conf_compute_rsci_biwt),
      .plm_conf_compute_rsci_bdwt(plm_conf_compute_rsci_bdwt),
      .plm_conf_compute_rsci_bcwt(plm_conf_compute_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci (
  clk, rst, plm_conf_load_rsc_dat, plm_conf_load_rsc_vld, plm_conf_load_rsc_rdy,
      core_wen, plm_conf_load_rsci_oswt_unreg, plm_conf_load_rsci_bawt, plm_conf_load_rsci_iswt0,
      plm_conf_load_rsci_wen_comp, plm_conf_load_rsci_idat
);
  input clk;
  input rst;
  output [255:0] plm_conf_load_rsc_dat;
  output plm_conf_load_rsc_vld;
  input plm_conf_load_rsc_rdy;
  input core_wen;
  input plm_conf_load_rsci_oswt_unreg;
  output plm_conf_load_rsci_bawt;
  input plm_conf_load_rsci_iswt0;
  output plm_conf_load_rsci_wen_comp;
  input [255:0] plm_conf_load_rsci_idat;


  // Interconnect Declarations
  wire plm_conf_load_rsci_irdy;
  wire plm_conf_load_rsci_biwt;
  wire plm_conf_load_rsci_bdwt;
  wire plm_conf_load_rsci_bcwt;
  wire plm_conf_load_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd256)) plm_conf_load_rsci (
      .irdy(plm_conf_load_rsci_irdy),
      .ivld(plm_conf_load_rsci_ivld_core_sct),
      .idat(plm_conf_load_rsci_idat),
      .rdy(plm_conf_load_rsc_rdy),
      .vld(plm_conf_load_rsc_vld),
      .dat(plm_conf_load_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl
      config_core_plm_conf_load_rsci_plm_conf_load_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_conf_load_rsci_oswt_unreg(plm_conf_load_rsci_oswt_unreg),
      .plm_conf_load_rsci_iswt0(plm_conf_load_rsci_iswt0),
      .plm_conf_load_rsci_irdy(plm_conf_load_rsci_irdy),
      .plm_conf_load_rsci_biwt(plm_conf_load_rsci_biwt),
      .plm_conf_load_rsci_bdwt(plm_conf_load_rsci_bdwt),
      .plm_conf_load_rsci_bcwt(plm_conf_load_rsci_bcwt),
      .plm_conf_load_rsci_ivld_core_sct(plm_conf_load_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci_plm_conf_load_wait_dp
      config_core_plm_conf_load_rsci_plm_conf_load_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_conf_load_rsci_oswt_unreg(plm_conf_load_rsci_oswt_unreg),
      .plm_conf_load_rsci_bawt(plm_conf_load_rsci_bawt),
      .plm_conf_load_rsci_wen_comp(plm_conf_load_rsci_wen_comp),
      .plm_conf_load_rsci_biwt(plm_conf_load_rsci_biwt),
      .plm_conf_load_rsci_bdwt(plm_conf_load_rsci_bdwt),
      .plm_conf_load_rsci_bcwt(plm_conf_load_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt_unreg,
      conf_info_rsci_bawt, conf_info_rsci_iswt0, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_wen_comp;
  output [255:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_ctrl config_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_iswt0(conf_info_rsci_iswt0),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci_conf_info_wait_dp config_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj (
  clk, rst, plm_filters_rsc_req_vz, core_wen, plm_filters_rsc_req_obj_oswt_unreg,
      plm_filters_rsc_req_obj_bawt, plm_filters_rsc_req_obj_iswt0, plm_filters_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_filters_rsc_req_vz;
  input core_wen;
  input plm_filters_rsc_req_obj_oswt_unreg;
  output plm_filters_rsc_req_obj_bawt;
  input plm_filters_rsc_req_obj_iswt0;
  output plm_filters_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_filters_rsc_req_obj_vd;
  wire plm_filters_rsc_req_obj_biwt;
  wire plm_filters_rsc_req_obj_bdwt;
  wire plm_filters_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_in_sync_v2 #(.valid(32'sd1)) plm_filters_rsc_req_obj
      (
      .vd(plm_filters_rsc_req_obj_vd),
      .vz(plm_filters_rsc_req_vz)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl
      load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_filters_rsc_req_obj_oswt_unreg(plm_filters_rsc_req_obj_oswt_unreg),
      .plm_filters_rsc_req_obj_iswt0(plm_filters_rsc_req_obj_iswt0),
      .plm_filters_rsc_req_obj_vd(plm_filters_rsc_req_obj_vd),
      .plm_filters_rsc_req_obj_biwt(plm_filters_rsc_req_obj_biwt),
      .plm_filters_rsc_req_obj_bdwt(plm_filters_rsc_req_obj_bdwt),
      .plm_filters_rsc_req_obj_bcwt(plm_filters_rsc_req_obj_bcwt)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp
      load_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_req_obj_oswt_unreg(plm_filters_rsc_req_obj_oswt_unreg),
      .plm_filters_rsc_req_obj_bawt(plm_filters_rsc_req_obj_bawt),
      .plm_filters_rsc_req_obj_wen_comp(plm_filters_rsc_req_obj_wen_comp),
      .plm_filters_rsc_req_obj_biwt(plm_filters_rsc_req_obj_biwt),
      .plm_filters_rsc_req_obj_bdwt(plm_filters_rsc_req_obj_bdwt),
      .plm_filters_rsc_req_obj_bcwt(plm_filters_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj (
  clk, rst, plm_inputs_rsc_req_vz, core_wen, plm_inputs_rsc_req_obj_oswt_unreg, plm_inputs_rsc_req_obj_bawt,
      plm_inputs_rsc_req_obj_iswt0, plm_inputs_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_inputs_rsc_req_vz;
  input core_wen;
  input plm_inputs_rsc_req_obj_oswt_unreg;
  output plm_inputs_rsc_req_obj_bawt;
  input plm_inputs_rsc_req_obj_iswt0;
  output plm_inputs_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_inputs_rsc_req_obj_vd;
  wire plm_inputs_rsc_req_obj_biwt;
  wire plm_inputs_rsc_req_obj_bdwt;
  wire plm_inputs_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_in_sync_v2 #(.valid(32'sd1)) plm_inputs_rsc_req_obj
      (
      .vd(plm_inputs_rsc_req_obj_vd),
      .vz(plm_inputs_rsc_req_vz)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl
      load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_inputs_rsc_req_obj_oswt_unreg(plm_inputs_rsc_req_obj_oswt_unreg),
      .plm_inputs_rsc_req_obj_iswt0(plm_inputs_rsc_req_obj_iswt0),
      .plm_inputs_rsc_req_obj_vd(plm_inputs_rsc_req_obj_vd),
      .plm_inputs_rsc_req_obj_biwt(plm_inputs_rsc_req_obj_biwt),
      .plm_inputs_rsc_req_obj_bdwt(plm_inputs_rsc_req_obj_bdwt),
      .plm_inputs_rsc_req_obj_bcwt(plm_inputs_rsc_req_obj_bcwt)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp
      load_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_req_obj_oswt_unreg(plm_inputs_rsc_req_obj_oswt_unreg),
      .plm_inputs_rsc_req_obj_bawt(plm_inputs_rsc_req_obj_bawt),
      .plm_inputs_rsc_req_obj_wen_comp(plm_inputs_rsc_req_obj_wen_comp),
      .plm_inputs_rsc_req_obj_biwt(plm_inputs_rsc_req_obj_biwt),
      .plm_inputs_rsc_req_obj_bdwt(plm_inputs_rsc_req_obj_bdwt),
      .plm_inputs_rsc_req_obj_bcwt(plm_inputs_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj (
  clk, rst, plm_filters_rsc_rls_lz, core_wen, core_wten, plm_filters_rsc_rls_obj_oswt_unreg,
      plm_filters_rsc_rls_obj_bawt, plm_filters_rsc_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_filters_rsc_rls_lz;
  input core_wen;
  input core_wten;
  input plm_filters_rsc_rls_obj_oswt_unreg;
  output plm_filters_rsc_rls_obj_bawt;
  input plm_filters_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_filters_rsc_rls_obj_biwt;
  wire plm_filters_rsc_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_io_sync_v2 #(.valid(32'sd0)) plm_filters_rsc_rls_obj
      (
      .ld(plm_filters_rsc_rls_obj_biwt),
      .lz(plm_filters_rsc_rls_lz)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl
      load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsc_rls_obj_oswt_unreg(plm_filters_rsc_rls_obj_oswt_unreg),
      .plm_filters_rsc_rls_obj_iswt0(plm_filters_rsc_rls_obj_iswt0),
      .plm_filters_rsc_rls_obj_biwt(plm_filters_rsc_rls_obj_biwt),
      .plm_filters_rsc_rls_obj_bdwt(plm_filters_rsc_rls_obj_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp
      load_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_rls_obj_bawt(plm_filters_rsc_rls_obj_bawt),
      .plm_filters_rsc_rls_obj_biwt(plm_filters_rsc_rls_obj_biwt),
      .plm_filters_rsc_rls_obj_bdwt(plm_filters_rsc_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj (
  clk, rst, plm_inputs_rsc_rls_lz, core_wen, core_wten, plm_inputs_rsc_rls_obj_oswt_unreg,
      plm_inputs_rsc_rls_obj_bawt, plm_inputs_rsc_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_inputs_rsc_rls_lz;
  input core_wen;
  input core_wten;
  input plm_inputs_rsc_rls_obj_oswt_unreg;
  output plm_inputs_rsc_rls_obj_bawt;
  input plm_inputs_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_inputs_rsc_rls_obj_biwt;
  wire plm_inputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_io_sync_v2 #(.valid(32'sd0)) plm_inputs_rsc_rls_obj
      (
      .ld(plm_inputs_rsc_rls_obj_biwt),
      .lz(plm_inputs_rsc_rls_lz)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl
      load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsc_rls_obj_oswt_unreg(plm_inputs_rsc_rls_obj_oswt_unreg),
      .plm_inputs_rsc_rls_obj_iswt0(plm_inputs_rsc_rls_obj_iswt0),
      .plm_inputs_rsc_rls_obj_biwt(plm_inputs_rsc_rls_obj_biwt),
      .plm_inputs_rsc_rls_obj_bdwt(plm_inputs_rsc_rls_obj_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp
      load_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_rls_obj_bawt(plm_inputs_rsc_rls_obj_bawt),
      .plm_inputs_rsc_rls_obj_biwt(plm_inputs_rsc_rls_obj_biwt),
      .plm_inputs_rsc_rls_obj_bdwt(plm_inputs_rsc_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt_unreg, done_rsci_bawt,
      done_rsci_iswt0, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  input done_rsci_iswt0;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd11)) done_rsci (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_load_core_done_rsci_done_wait_ctrl load_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_iswt0(done_rsci_iswt0),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_load_core_done_rsci_done_wait_dp load_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci (
  clk, rst, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy,
      core_wen, dma_read_chnl_rsci_oswt_unreg, dma_read_chnl_rsci_bawt, dma_read_chnl_rsci_iswt0,
      dma_read_chnl_rsci_wen_comp, dma_read_chnl_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  input core_wen;
  input dma_read_chnl_rsci_oswt_unreg;
  output dma_read_chnl_rsci_bawt;
  input dma_read_chnl_rsci_iswt0;
  output dma_read_chnl_rsci_wen_comp;
  output [31:0] dma_read_chnl_rsci_idat_mxwt;


  // Interconnect Declarations
  wire dma_read_chnl_rsci_biwt;
  wire dma_read_chnl_rsci_bdwt;
  wire dma_read_chnl_rsci_bcwt;
  wire dma_read_chnl_rsci_irdy_core_sct;
  wire dma_read_chnl_rsci_ivld;
  wire [63:0] dma_read_chnl_rsci_idat;
  wire [31:0] dma_read_chnl_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd10),
  .width(32'sd64)) dma_read_chnl_rsci (
      .rdy(dma_read_chnl_rsc_rdy),
      .vld(dma_read_chnl_rsc_vld),
      .dat(dma_read_chnl_rsc_dat),
      .irdy(dma_read_chnl_rsci_irdy_core_sct),
      .ivld(dma_read_chnl_rsci_ivld),
      .idat(dma_read_chnl_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl
      load_core_dma_read_chnl_rsci_dma_read_chnl_wait_ctrl_inst (
      .core_wen(core_wen),
      .dma_read_chnl_rsci_oswt_unreg(dma_read_chnl_rsci_oswt_unreg),
      .dma_read_chnl_rsci_iswt0(dma_read_chnl_rsci_iswt0),
      .dma_read_chnl_rsci_biwt(dma_read_chnl_rsci_biwt),
      .dma_read_chnl_rsci_bdwt(dma_read_chnl_rsci_bdwt),
      .dma_read_chnl_rsci_bcwt(dma_read_chnl_rsci_bcwt),
      .dma_read_chnl_rsci_irdy_core_sct(dma_read_chnl_rsci_irdy_core_sct),
      .dma_read_chnl_rsci_ivld(dma_read_chnl_rsci_ivld)
    );
  esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp
      load_core_dma_read_chnl_rsci_dma_read_chnl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_rsci_oswt_unreg(dma_read_chnl_rsci_oswt_unreg),
      .dma_read_chnl_rsci_bawt(dma_read_chnl_rsci_bawt),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .dma_read_chnl_rsci_idat_mxwt(dma_read_chnl_rsci_idat_mxwt_pconst),
      .dma_read_chnl_rsci_biwt(dma_read_chnl_rsci_biwt),
      .dma_read_chnl_rsci_bdwt(dma_read_chnl_rsci_bdwt),
      .dma_read_chnl_rsci_bcwt(dma_read_chnl_rsci_bcwt),
      .dma_read_chnl_rsci_idat(dma_read_chnl_rsci_idat)
    );
  assign dma_read_chnl_rsci_idat_mxwt = dma_read_chnl_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci (
  clk, rst, dma_read_ctrl_rsc_dat, dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy,
      core_wen, core_wten, dma_read_ctrl_rsci_oswt_unreg, dma_read_ctrl_rsci_bawt,
      dma_read_ctrl_rsci_iswt0, dma_read_ctrl_rsci_irdy_mxwt, dma_read_ctrl_rsci_idat
);
  input clk;
  input rst;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  input core_wen;
  input core_wten;
  input dma_read_ctrl_rsci_oswt_unreg;
  output dma_read_ctrl_rsci_bawt;
  input dma_read_ctrl_rsci_iswt0;
  output dma_read_ctrl_rsci_irdy_mxwt;
  input [66:0] dma_read_ctrl_rsci_idat;


  // Interconnect Declarations
  wire dma_read_ctrl_rsci_irdy;
  wire dma_read_ctrl_rsci_biwt;
  wire dma_read_ctrl_rsci_bdwt;


  // Interconnect Declarations for Component Instantiations 
  wire [66:0] nl_dma_read_ctrl_rsci_idat;
  assign nl_dma_read_ctrl_rsci_idat = {19'b0110000000000000000 , (dma_read_ctrl_rsci_idat[47:32])
      , 16'b0000000000000000 , (dma_read_ctrl_rsci_idat[15:0])};
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd9),
  .width(32'sd67)) dma_read_ctrl_rsci (
      .irdy(dma_read_ctrl_rsci_irdy),
      .ivld(dma_read_ctrl_rsci_biwt),
      .idat(nl_dma_read_ctrl_rsci_idat[66:0]),
      .rdy(dma_read_ctrl_rsc_rdy),
      .vld(dma_read_ctrl_rsc_vld),
      .dat(dma_read_ctrl_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl
      load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dma_read_ctrl_rsci_oswt_unreg(dma_read_ctrl_rsci_oswt_unreg),
      .dma_read_ctrl_rsci_iswt0(dma_read_ctrl_rsci_iswt0),
      .dma_read_ctrl_rsci_biwt(dma_read_ctrl_rsci_biwt),
      .dma_read_ctrl_rsci_bdwt(dma_read_ctrl_rsci_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp
      load_core_dma_read_ctrl_rsci_dma_read_ctrl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_rsci_bawt(dma_read_ctrl_rsci_bawt),
      .dma_read_ctrl_rsci_irdy_mxwt(dma_read_ctrl_rsci_irdy_mxwt),
      .dma_read_ctrl_rsci_irdy(dma_read_ctrl_rsci_irdy),
      .dma_read_ctrl_rsci_biwt(dma_read_ctrl_rsci_biwt),
      .dma_read_ctrl_rsci_bdwt(dma_read_ctrl_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1 (
  clk, rst, core_wen, core_wten, plm_filters_rsci_oswt_unreg, plm_filters_rsci_bawt,
      plm_filters_rsci_iswt0, plm_filters_rsci_we_d_pff, plm_filters_rsci_iswt0_pff
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input plm_filters_rsci_oswt_unreg;
  output plm_filters_rsci_bawt;
  input plm_filters_rsci_iswt0;
  output plm_filters_rsci_we_d_pff;
  input plm_filters_rsci_iswt0_pff;


  // Interconnect Declarations
  wire plm_filters_rsci_biwt;
  wire plm_filters_rsci_bdwt;
  wire plm_filters_rsci_we_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl
      load_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsci_oswt_unreg(plm_filters_rsci_oswt_unreg),
      .plm_filters_rsci_iswt0(plm_filters_rsci_iswt0),
      .plm_filters_rsci_biwt(plm_filters_rsci_biwt),
      .plm_filters_rsci_bdwt(plm_filters_rsci_bdwt),
      .plm_filters_rsci_we_d_core_sct_pff(plm_filters_rsci_we_d_core_sct_iff),
      .plm_filters_rsci_iswt0_pff(plm_filters_rsci_iswt0_pff)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp
      load_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsci_bawt(plm_filters_rsci_bawt),
      .plm_filters_rsci_biwt(plm_filters_rsci_biwt),
      .plm_filters_rsci_bdwt(plm_filters_rsci_bdwt)
    );
  assign plm_filters_rsci_we_d_pff = plm_filters_rsci_we_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1 (
  clk, rst, core_wen, core_wten, plm_inputs_rsci_oswt_unreg, plm_inputs_rsci_bawt,
      plm_inputs_rsci_iswt0, plm_inputs_rsci_we_d_pff, plm_inputs_rsci_iswt0_pff
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input plm_inputs_rsci_oswt_unreg;
  output plm_inputs_rsci_bawt;
  input plm_inputs_rsci_iswt0;
  output plm_inputs_rsci_we_d_pff;
  input plm_inputs_rsci_iswt0_pff;


  // Interconnect Declarations
  wire plm_inputs_rsci_biwt;
  wire plm_inputs_rsci_bdwt;
  wire plm_inputs_rsci_we_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl
      load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsci_oswt_unreg(plm_inputs_rsci_oswt_unreg),
      .plm_inputs_rsci_iswt0(plm_inputs_rsci_iswt0),
      .plm_inputs_rsci_biwt(plm_inputs_rsci_biwt),
      .plm_inputs_rsci_bdwt(plm_inputs_rsci_bdwt),
      .plm_inputs_rsci_we_d_core_sct_pff(plm_inputs_rsci_we_d_core_sct_iff),
      .plm_inputs_rsci_iswt0_pff(plm_inputs_rsci_iswt0_pff)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp
      load_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsci_bawt(plm_inputs_rsci_bawt),
      .plm_inputs_rsci_biwt(plm_inputs_rsci_biwt),
      .plm_inputs_rsci_bdwt(plm_inputs_rsci_bdwt)
    );
  assign plm_inputs_rsci_we_d_pff = plm_inputs_rsci_we_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt_unreg,
      conf_info_rsci_bawt, conf_info_rsci_iswt0, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;
  wire [63:0] conf_info_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd6),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_ctrl load_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_iswt0(conf_info_rsci_iswt0),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci_conf_info_wait_dp load_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt_pconst),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
  assign conf_info_rsci_idat_mxwt = conf_info_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj (
  clk, rst, plm_outputs_rsc_req_vz, core_wen, plm_outputs_rsc_req_obj_oswt_unreg,
      plm_outputs_rsc_req_obj_bawt, plm_outputs_rsc_req_obj_iswt0, plm_outputs_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_outputs_rsc_req_vz;
  input core_wen;
  input plm_outputs_rsc_req_obj_oswt_unreg;
  output plm_outputs_rsc_req_obj_bawt;
  input plm_outputs_rsc_req_obj_iswt0;
  output plm_outputs_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_outputs_rsc_req_obj_vd;
  wire plm_outputs_rsc_req_obj_biwt;
  wire plm_outputs_rsc_req_obj_bdwt;
  wire plm_outputs_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_in_sync_v2 #(.valid(32'sd1)) plm_outputs_rsc_req_obj
      (
      .vd(plm_outputs_rsc_req_obj_vd),
      .vz(plm_outputs_rsc_req_vz)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl
      compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_outputs_rsc_req_obj_oswt_unreg(plm_outputs_rsc_req_obj_oswt_unreg),
      .plm_outputs_rsc_req_obj_iswt0(plm_outputs_rsc_req_obj_iswt0),
      .plm_outputs_rsc_req_obj_vd(plm_outputs_rsc_req_obj_vd),
      .plm_outputs_rsc_req_obj_biwt(plm_outputs_rsc_req_obj_biwt),
      .plm_outputs_rsc_req_obj_bdwt(plm_outputs_rsc_req_obj_bdwt),
      .plm_outputs_rsc_req_obj_bcwt(plm_outputs_rsc_req_obj_bcwt)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp
      compute_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_req_obj_oswt_unreg(plm_outputs_rsc_req_obj_oswt_unreg),
      .plm_outputs_rsc_req_obj_bawt(plm_outputs_rsc_req_obj_bawt),
      .plm_outputs_rsc_req_obj_wen_comp(plm_outputs_rsc_req_obj_wen_comp),
      .plm_outputs_rsc_req_obj_biwt(plm_outputs_rsc_req_obj_biwt),
      .plm_outputs_rsc_req_obj_bdwt(plm_outputs_rsc_req_obj_bdwt),
      .plm_outputs_rsc_req_obj_bcwt(plm_outputs_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj (
  clk, rst, plm_inputs_rsc_req_vz, core_wen, plm_inputs_rsc_req_obj_oswt_unreg, plm_inputs_rsc_req_obj_bawt,
      plm_inputs_rsc_req_obj_iswt0, plm_inputs_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_inputs_rsc_req_vz;
  input core_wen;
  input plm_inputs_rsc_req_obj_oswt_unreg;
  output plm_inputs_rsc_req_obj_bawt;
  input plm_inputs_rsc_req_obj_iswt0;
  output plm_inputs_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_inputs_rsc_req_obj_vd;
  wire plm_inputs_rsc_req_obj_biwt;
  wire plm_inputs_rsc_req_obj_bdwt;
  wire plm_inputs_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_in_sync_v2 #(.valid(32'sd1)) plm_inputs_rsc_req_obj
      (
      .vd(plm_inputs_rsc_req_obj_vd),
      .vz(plm_inputs_rsc_req_vz)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl
      compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_inputs_rsc_req_obj_oswt_unreg(plm_inputs_rsc_req_obj_oswt_unreg),
      .plm_inputs_rsc_req_obj_iswt0(plm_inputs_rsc_req_obj_iswt0),
      .plm_inputs_rsc_req_obj_vd(plm_inputs_rsc_req_obj_vd),
      .plm_inputs_rsc_req_obj_biwt(plm_inputs_rsc_req_obj_biwt),
      .plm_inputs_rsc_req_obj_bdwt(plm_inputs_rsc_req_obj_bdwt),
      .plm_inputs_rsc_req_obj_bcwt(plm_inputs_rsc_req_obj_bcwt)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp
      compute_core_plm_inputs_rsc_req_obj_plm_inputs_rsc_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_req_obj_oswt_unreg(plm_inputs_rsc_req_obj_oswt_unreg),
      .plm_inputs_rsc_req_obj_bawt(plm_inputs_rsc_req_obj_bawt),
      .plm_inputs_rsc_req_obj_wen_comp(plm_inputs_rsc_req_obj_wen_comp),
      .plm_inputs_rsc_req_obj_biwt(plm_inputs_rsc_req_obj_biwt),
      .plm_inputs_rsc_req_obj_bdwt(plm_inputs_rsc_req_obj_bdwt),
      .plm_inputs_rsc_req_obj_bcwt(plm_inputs_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj (
  clk, rst, plm_filters_rsc_req_vz, core_wen, plm_filters_rsc_req_obj_oswt_unreg,
      plm_filters_rsc_req_obj_bawt, plm_filters_rsc_req_obj_iswt0, plm_filters_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_filters_rsc_req_vz;
  input core_wen;
  input plm_filters_rsc_req_obj_oswt_unreg;
  output plm_filters_rsc_req_obj_bawt;
  input plm_filters_rsc_req_obj_iswt0;
  output plm_filters_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_filters_rsc_req_obj_vd;
  wire plm_filters_rsc_req_obj_biwt;
  wire plm_filters_rsc_req_obj_bdwt;
  wire plm_filters_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_in_sync_v2 #(.valid(32'sd1)) plm_filters_rsc_req_obj
      (
      .vd(plm_filters_rsc_req_obj_vd),
      .vz(plm_filters_rsc_req_vz)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl
      compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_filters_rsc_req_obj_oswt_unreg(plm_filters_rsc_req_obj_oswt_unreg),
      .plm_filters_rsc_req_obj_iswt0(plm_filters_rsc_req_obj_iswt0),
      .plm_filters_rsc_req_obj_vd(plm_filters_rsc_req_obj_vd),
      .plm_filters_rsc_req_obj_biwt(plm_filters_rsc_req_obj_biwt),
      .plm_filters_rsc_req_obj_bdwt(plm_filters_rsc_req_obj_bdwt),
      .plm_filters_rsc_req_obj_bcwt(plm_filters_rsc_req_obj_bcwt)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp
      compute_core_plm_filters_rsc_req_obj_plm_filters_rsc_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_req_obj_oswt_unreg(plm_filters_rsc_req_obj_oswt_unreg),
      .plm_filters_rsc_req_obj_bawt(plm_filters_rsc_req_obj_bawt),
      .plm_filters_rsc_req_obj_wen_comp(plm_filters_rsc_req_obj_wen_comp),
      .plm_filters_rsc_req_obj_biwt(plm_filters_rsc_req_obj_biwt),
      .plm_filters_rsc_req_obj_bdwt(plm_filters_rsc_req_obj_bdwt),
      .plm_filters_rsc_req_obj_bcwt(plm_filters_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj (
  clk, rst, plm_filters_rsc_rls_lz, core_wen, core_wten, plm_filters_rsc_rls_obj_oswt_unreg,
      plm_filters_rsc_rls_obj_bawt, plm_filters_rsc_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_filters_rsc_rls_lz;
  input core_wen;
  input core_wten;
  input plm_filters_rsc_rls_obj_oswt_unreg;
  output plm_filters_rsc_rls_obj_bawt;
  input plm_filters_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_filters_rsc_rls_obj_biwt;
  wire plm_filters_rsc_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_io_sync_v2 #(.valid(32'sd0)) plm_filters_rsc_rls_obj
      (
      .ld(plm_filters_rsc_rls_obj_biwt),
      .lz(plm_filters_rsc_rls_lz)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl
      compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsc_rls_obj_oswt_unreg(plm_filters_rsc_rls_obj_oswt_unreg),
      .plm_filters_rsc_rls_obj_iswt0(plm_filters_rsc_rls_obj_iswt0),
      .plm_filters_rsc_rls_obj_biwt(plm_filters_rsc_rls_obj_biwt),
      .plm_filters_rsc_rls_obj_bdwt(plm_filters_rsc_rls_obj_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp
      compute_core_plm_filters_rsc_rls_obj_plm_filters_rsc_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_rls_obj_bawt(plm_filters_rsc_rls_obj_bawt),
      .plm_filters_rsc_rls_obj_biwt(plm_filters_rsc_rls_obj_biwt),
      .plm_filters_rsc_rls_obj_bdwt(plm_filters_rsc_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj (
  clk, rst, plm_inputs_rsc_rls_lz, core_wen, core_wten, plm_inputs_rsc_rls_obj_oswt_unreg,
      plm_inputs_rsc_rls_obj_bawt, plm_inputs_rsc_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_inputs_rsc_rls_lz;
  input core_wen;
  input core_wten;
  input plm_inputs_rsc_rls_obj_oswt_unreg;
  output plm_inputs_rsc_rls_obj_bawt;
  input plm_inputs_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_inputs_rsc_rls_obj_biwt;
  wire plm_inputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_io_sync_v2 #(.valid(32'sd0)) plm_inputs_rsc_rls_obj
      (
      .ld(plm_inputs_rsc_rls_obj_biwt),
      .lz(plm_inputs_rsc_rls_lz)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl
      compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsc_rls_obj_oswt_unreg(plm_inputs_rsc_rls_obj_oswt_unreg),
      .plm_inputs_rsc_rls_obj_iswt0(plm_inputs_rsc_rls_obj_iswt0),
      .plm_inputs_rsc_rls_obj_biwt(plm_inputs_rsc_rls_obj_biwt),
      .plm_inputs_rsc_rls_obj_bdwt(plm_inputs_rsc_rls_obj_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp
      compute_core_plm_inputs_rsc_rls_obj_plm_inputs_rsc_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_rls_obj_bawt(plm_inputs_rsc_rls_obj_bawt),
      .plm_inputs_rsc_rls_obj_biwt(plm_inputs_rsc_rls_obj_biwt),
      .plm_inputs_rsc_rls_obj_bdwt(plm_inputs_rsc_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj (
  clk, rst, plm_outputs_rsc_rls_lz, core_wen, core_wten, plm_outputs_rsc_rls_obj_oswt_unreg,
      plm_outputs_rsc_rls_obj_bawt, plm_outputs_rsc_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_outputs_rsc_rls_lz;
  input core_wen;
  input core_wten;
  input plm_outputs_rsc_rls_obj_oswt_unreg;
  output plm_outputs_rsc_rls_obj_bawt;
  input plm_outputs_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_outputs_rsc_rls_obj_biwt;
  wire plm_outputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_io_sync_v2 #(.valid(32'sd0)) plm_outputs_rsc_rls_obj
      (
      .ld(plm_outputs_rsc_rls_obj_biwt),
      .lz(plm_outputs_rsc_rls_lz)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl
      compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsc_rls_obj_oswt_unreg(plm_outputs_rsc_rls_obj_oswt_unreg),
      .plm_outputs_rsc_rls_obj_iswt0(plm_outputs_rsc_rls_obj_iswt0),
      .plm_outputs_rsc_rls_obj_biwt(plm_outputs_rsc_rls_obj_biwt),
      .plm_outputs_rsc_rls_obj_bdwt(plm_outputs_rsc_rls_obj_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp
      compute_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_rls_obj_bawt(plm_outputs_rsc_rls_obj_bawt),
      .plm_outputs_rsc_rls_obj_biwt(plm_outputs_rsc_rls_obj_biwt),
      .plm_outputs_rsc_rls_obj_bdwt(plm_outputs_rsc_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt_unreg, done_rsci_bawt,
      done_rsci_iswt0, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  input done_rsci_iswt0;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd18)) done_rsci (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_done_rsci_done_wait_ctrl compute_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_iswt0(done_rsci_iswt0),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_done_rsci_done_wait_dp compute_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1 (
  clk, rst, core_wen, core_wten, plm_outputs_rsci_oswt_unreg, plm_outputs_rsci_bawt,
      plm_outputs_rsci_iswt0, plm_outputs_rsci_we_d_pff, plm_outputs_rsci_iswt0_pff
);
  input clk;
  input rst;
  input core_wen;
  input core_wten;
  input plm_outputs_rsci_oswt_unreg;
  output plm_outputs_rsci_bawt;
  input plm_outputs_rsci_iswt0;
  output plm_outputs_rsci_we_d_pff;
  input plm_outputs_rsci_iswt0_pff;


  // Interconnect Declarations
  wire plm_outputs_rsci_biwt;
  wire plm_outputs_rsci_bdwt;
  wire plm_outputs_rsci_we_d_core_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl
      compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsci_oswt_unreg(plm_outputs_rsci_oswt_unreg),
      .plm_outputs_rsci_iswt0(plm_outputs_rsci_iswt0),
      .plm_outputs_rsci_biwt(plm_outputs_rsci_biwt),
      .plm_outputs_rsci_bdwt(plm_outputs_rsci_bdwt),
      .plm_outputs_rsci_we_d_core_sct_pff(plm_outputs_rsci_we_d_core_sct_iff),
      .plm_outputs_rsci_iswt0_pff(plm_outputs_rsci_iswt0_pff)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp
      compute_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsci_bawt(plm_outputs_rsci_bawt),
      .plm_outputs_rsci_biwt(plm_outputs_rsci_biwt),
      .plm_outputs_rsci_bdwt(plm_outputs_rsci_bdwt)
    );
  assign plm_outputs_rsci_we_d_pff = plm_outputs_rsci_we_d_core_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1 (
  clk, rst, plm_filters_rsci_q_d, plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, plm_filters_rsci_oswt_unreg, plm_filters_rsci_bawt, plm_filters_rsci_iswt0,
      plm_filters_rsci_q_d_mxwt, plm_filters_rsci_iswt0_pff
);
  input clk;
  input rst;
  input [31:0] plm_filters_rsci_q_d;
  output plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input plm_filters_rsci_oswt_unreg;
  output plm_filters_rsci_bawt;
  input plm_filters_rsci_iswt0;
  output [31:0] plm_filters_rsci_q_d_mxwt;
  input plm_filters_rsci_iswt0_pff;


  // Interconnect Declarations
  wire plm_filters_rsci_biwt;
  wire plm_filters_rsci_bdwt;
  wire plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl
      compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsci_oswt_unreg(plm_filters_rsci_oswt_unreg),
      .plm_filters_rsci_iswt0(plm_filters_rsci_iswt0),
      .plm_filters_rsci_biwt(plm_filters_rsci_biwt),
      .plm_filters_rsci_bdwt(plm_filters_rsci_bdwt),
      .plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct(plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct),
      .plm_filters_rsci_iswt0_pff(plm_filters_rsci_iswt0_pff)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp
      compute_core_plm_filters_rsci_1_plm_filters_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsci_q_d(plm_filters_rsci_q_d),
      .plm_filters_rsci_bawt(plm_filters_rsci_bawt),
      .plm_filters_rsci_q_d_mxwt(plm_filters_rsci_q_d_mxwt),
      .plm_filters_rsci_biwt(plm_filters_rsci_biwt),
      .plm_filters_rsci_bdwt(plm_filters_rsci_bdwt)
    );
  assign plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1 (
  clk, rst, plm_inputs_rsci_q_d, plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, plm_inputs_rsci_oswt_unreg, plm_inputs_rsci_bawt, plm_inputs_rsci_iswt0,
      plm_inputs_rsci_q_d_mxwt, plm_inputs_rsci_iswt0_pff
);
  input clk;
  input rst;
  input [31:0] plm_inputs_rsci_q_d;
  output plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input plm_inputs_rsci_oswt_unreg;
  output plm_inputs_rsci_bawt;
  input plm_inputs_rsci_iswt0;
  output [31:0] plm_inputs_rsci_q_d_mxwt;
  input plm_inputs_rsci_iswt0_pff;


  // Interconnect Declarations
  wire plm_inputs_rsci_biwt;
  wire plm_inputs_rsci_bdwt;
  wire plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl
      compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsci_oswt_unreg(plm_inputs_rsci_oswt_unreg),
      .plm_inputs_rsci_iswt0(plm_inputs_rsci_iswt0),
      .plm_inputs_rsci_biwt(plm_inputs_rsci_biwt),
      .plm_inputs_rsci_bdwt(plm_inputs_rsci_bdwt),
      .plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct(plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct),
      .plm_inputs_rsci_iswt0_pff(plm_inputs_rsci_iswt0_pff)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp
      compute_core_plm_inputs_rsci_1_plm_inputs_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsci_q_d(plm_inputs_rsci_q_d),
      .plm_inputs_rsci_bawt(plm_inputs_rsci_bawt),
      .plm_inputs_rsci_q_d_mxwt(plm_inputs_rsci_q_d_mxwt),
      .plm_inputs_rsci_biwt(plm_inputs_rsci_biwt),
      .plm_inputs_rsci_bdwt(plm_inputs_rsci_bdwt)
    );
  assign plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt_unreg,
      conf_info_rsci_bawt, conf_info_rsci_iswt0, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;
  wire [63:0] conf_info_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd14),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_ctrl compute_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_iswt0(conf_info_rsci_iswt0),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci_conf_info_wait_dp compute_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt_pconst),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
  assign conf_info_rsci_idat_mxwt = conf_info_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj (
  clk, rst, plm_outputs_rsc_req_vz, core_wen, plm_outputs_rsc_req_obj_oswt_unreg,
      plm_outputs_rsc_req_obj_bawt, plm_outputs_rsc_req_obj_iswt0, plm_outputs_rsc_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_outputs_rsc_req_vz;
  input core_wen;
  input plm_outputs_rsc_req_obj_oswt_unreg;
  output plm_outputs_rsc_req_obj_bawt;
  input plm_outputs_rsc_req_obj_iswt0;
  output plm_outputs_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_outputs_rsc_req_obj_vd;
  wire plm_outputs_rsc_req_obj_biwt;
  wire plm_outputs_rsc_req_obj_bdwt;
  wire plm_outputs_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_in_sync_v2 #(.valid(32'sd1)) plm_outputs_rsc_req_obj
      (
      .vd(plm_outputs_rsc_req_obj_vd),
      .vz(plm_outputs_rsc_req_vz)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl
      store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_ctrl_inst (
      .core_wen(core_wen),
      .plm_outputs_rsc_req_obj_oswt_unreg(plm_outputs_rsc_req_obj_oswt_unreg),
      .plm_outputs_rsc_req_obj_iswt0(plm_outputs_rsc_req_obj_iswt0),
      .plm_outputs_rsc_req_obj_vd(plm_outputs_rsc_req_obj_vd),
      .plm_outputs_rsc_req_obj_biwt(plm_outputs_rsc_req_obj_biwt),
      .plm_outputs_rsc_req_obj_bdwt(plm_outputs_rsc_req_obj_bdwt),
      .plm_outputs_rsc_req_obj_bcwt(plm_outputs_rsc_req_obj_bcwt)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp
      store_core_plm_outputs_rsc_req_obj_plm_outputs_rsc_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_req_obj_oswt_unreg(plm_outputs_rsc_req_obj_oswt_unreg),
      .plm_outputs_rsc_req_obj_bawt(plm_outputs_rsc_req_obj_bawt),
      .plm_outputs_rsc_req_obj_wen_comp(plm_outputs_rsc_req_obj_wen_comp),
      .plm_outputs_rsc_req_obj_biwt(plm_outputs_rsc_req_obj_biwt),
      .plm_outputs_rsc_req_obj_bdwt(plm_outputs_rsc_req_obj_bdwt),
      .plm_outputs_rsc_req_obj_bcwt(plm_outputs_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj (
  clk, rst, plm_outputs_rsc_rls_lz, core_wen, core_wten, plm_outputs_rsc_rls_obj_oswt_unreg,
      plm_outputs_rsc_rls_obj_bawt, plm_outputs_rsc_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_outputs_rsc_rls_lz;
  input core_wen;
  input core_wten;
  input plm_outputs_rsc_rls_obj_oswt_unreg;
  output plm_outputs_rsc_rls_obj_bawt;
  input plm_outputs_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_outputs_rsc_rls_obj_biwt;
  wire plm_outputs_rsc_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_mgc_io_sync_v2 #(.valid(32'sd0)) plm_outputs_rsc_rls_obj
      (
      .ld(plm_outputs_rsc_rls_obj_biwt),
      .lz(plm_outputs_rsc_rls_lz)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl
      store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsc_rls_obj_oswt_unreg(plm_outputs_rsc_rls_obj_oswt_unreg),
      .plm_outputs_rsc_rls_obj_iswt0(plm_outputs_rsc_rls_obj_iswt0),
      .plm_outputs_rsc_rls_obj_biwt(plm_outputs_rsc_rls_obj_biwt),
      .plm_outputs_rsc_rls_obj_bdwt(plm_outputs_rsc_rls_obj_bdwt)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp
      store_core_plm_outputs_rsc_rls_obj_plm_outputs_rsc_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_rls_obj_bawt(plm_outputs_rsc_rls_obj_bawt),
      .plm_outputs_rsc_rls_obj_biwt(plm_outputs_rsc_rls_obj_biwt),
      .plm_outputs_rsc_rls_obj_bdwt(plm_outputs_rsc_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_done_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_done_rsci (
  clk, rst, done_rsc_rdy, done_rsc_vld, core_wen, done_rsci_oswt_unreg, done_rsci_bawt,
      done_rsci_iswt0, done_rsci_wen_comp
);
  input clk;
  input rst;
  input done_rsc_rdy;
  output done_rsc_vld;
  input core_wen;
  input done_rsci_oswt_unreg;
  output done_rsci_bawt;
  input done_rsci_iswt0;
  output done_rsci_wen_comp;


  // Interconnect Declarations
  wire done_rsci_biwt;
  wire done_rsci_bdwt;
  wire done_rsci_bcwt;
  wire done_rsci_ivld_core_sct;
  wire done_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_sync_out_wait_v1 #(.rscid(32'sd27)) done_rsci (
      .vld(done_rsc_vld),
      .rdy(done_rsc_rdy),
      .ivld(done_rsci_ivld_core_sct),
      .irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_store_core_done_rsci_done_wait_ctrl store_core_done_rsci_done_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_iswt0(done_rsci_iswt0),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt),
      .done_rsci_ivld_core_sct(done_rsci_ivld_core_sct),
      .done_rsci_irdy(done_rsci_irdy)
    );
  esp_acc_conv2d_cxx_catapult_store_core_done_rsci_done_wait_dp store_core_done_rsci_done_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsci_oswt_unreg(done_rsci_oswt_unreg),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .done_rsci_biwt(done_rsci_biwt),
      .done_rsci_bdwt(done_rsci_bdwt),
      .done_rsci_bcwt(done_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci (
  clk, rst, dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy,
      core_wen, dma_write_chnl_rsci_oswt_unreg, dma_write_chnl_rsci_bawt, dma_write_chnl_rsci_iswt0,
      dma_write_chnl_rsci_wen_comp, dma_write_chnl_rsci_idat
);
  input clk;
  input rst;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  input core_wen;
  input dma_write_chnl_rsci_oswt_unreg;
  output dma_write_chnl_rsci_bawt;
  input dma_write_chnl_rsci_iswt0;
  output dma_write_chnl_rsci_wen_comp;
  input [63:0] dma_write_chnl_rsci_idat;


  // Interconnect Declarations
  wire dma_write_chnl_rsci_irdy;
  wire dma_write_chnl_rsci_biwt;
  wire dma_write_chnl_rsci_bdwt;
  wire dma_write_chnl_rsci_bcwt;
  wire dma_write_chnl_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_dma_write_chnl_rsci_idat;
  assign nl_dma_write_chnl_rsci_idat = {32'b11011110101011011011111011101111 , (dma_write_chnl_rsci_idat[31:0])};
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd26),
  .width(32'sd64)) dma_write_chnl_rsci (
      .irdy(dma_write_chnl_rsci_irdy),
      .ivld(dma_write_chnl_rsci_ivld_core_sct),
      .idat(nl_dma_write_chnl_rsci_idat[63:0]),
      .rdy(dma_write_chnl_rsc_rdy),
      .vld(dma_write_chnl_rsc_vld),
      .dat(dma_write_chnl_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl
      store_core_dma_write_chnl_rsci_dma_write_chnl_wait_ctrl_inst (
      .core_wen(core_wen),
      .dma_write_chnl_rsci_oswt_unreg(dma_write_chnl_rsci_oswt_unreg),
      .dma_write_chnl_rsci_iswt0(dma_write_chnl_rsci_iswt0),
      .dma_write_chnl_rsci_irdy(dma_write_chnl_rsci_irdy),
      .dma_write_chnl_rsci_biwt(dma_write_chnl_rsci_biwt),
      .dma_write_chnl_rsci_bdwt(dma_write_chnl_rsci_bdwt),
      .dma_write_chnl_rsci_bcwt(dma_write_chnl_rsci_bcwt),
      .dma_write_chnl_rsci_ivld_core_sct(dma_write_chnl_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp
      store_core_dma_write_chnl_rsci_dma_write_chnl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_rsci_oswt_unreg(dma_write_chnl_rsci_oswt_unreg),
      .dma_write_chnl_rsci_bawt(dma_write_chnl_rsci_bawt),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .dma_write_chnl_rsci_biwt(dma_write_chnl_rsci_biwt),
      .dma_write_chnl_rsci_bdwt(dma_write_chnl_rsci_bdwt),
      .dma_write_chnl_rsci_bcwt(dma_write_chnl_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci (
  clk, rst, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy,
      core_wen, dma_write_ctrl_rsci_oswt_unreg, dma_write_ctrl_rsci_bawt, dma_write_ctrl_rsci_iswt0,
      dma_write_ctrl_rsci_wen_comp, dma_write_ctrl_rsci_idat
);
  input clk;
  input rst;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input core_wen;
  input dma_write_ctrl_rsci_oswt_unreg;
  output dma_write_ctrl_rsci_bawt;
  input dma_write_ctrl_rsci_iswt0;
  output dma_write_ctrl_rsci_wen_comp;
  input [66:0] dma_write_ctrl_rsci_idat;


  // Interconnect Declarations
  wire dma_write_ctrl_rsci_irdy;
  wire dma_write_ctrl_rsci_biwt;
  wire dma_write_ctrl_rsci_bdwt;
  wire dma_write_ctrl_rsci_bcwt;
  wire dma_write_ctrl_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [66:0] nl_dma_write_ctrl_rsci_idat;
  assign nl_dma_write_ctrl_rsci_idat = {19'b0110000000000000000 , (dma_write_ctrl_rsci_idat[47:32])
      , 16'b0000000000000000 , (dma_write_ctrl_rsci_idat[15:0])};
  esp_acc_conv2d_cxx_catapult_ccs_out_wait_v1 #(.rscid(32'sd25),
  .width(32'sd67)) dma_write_ctrl_rsci (
      .irdy(dma_write_ctrl_rsci_irdy),
      .ivld(dma_write_ctrl_rsci_ivld_core_sct),
      .idat(nl_dma_write_ctrl_rsci_idat[66:0]),
      .rdy(dma_write_ctrl_rsc_rdy),
      .vld(dma_write_ctrl_rsc_vld),
      .dat(dma_write_ctrl_rsc_dat)
    );
  esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl
      store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_ctrl_inst (
      .core_wen(core_wen),
      .dma_write_ctrl_rsci_oswt_unreg(dma_write_ctrl_rsci_oswt_unreg),
      .dma_write_ctrl_rsci_iswt0(dma_write_ctrl_rsci_iswt0),
      .dma_write_ctrl_rsci_irdy(dma_write_ctrl_rsci_irdy),
      .dma_write_ctrl_rsci_biwt(dma_write_ctrl_rsci_biwt),
      .dma_write_ctrl_rsci_bdwt(dma_write_ctrl_rsci_bdwt),
      .dma_write_ctrl_rsci_bcwt(dma_write_ctrl_rsci_bcwt),
      .dma_write_ctrl_rsci_ivld_core_sct(dma_write_ctrl_rsci_ivld_core_sct)
    );
  esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp
      store_core_dma_write_ctrl_rsci_dma_write_ctrl_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_rsci_oswt_unreg(dma_write_ctrl_rsci_oswt_unreg),
      .dma_write_ctrl_rsci_bawt(dma_write_ctrl_rsci_bawt),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_ctrl_rsci_biwt(dma_write_ctrl_rsci_biwt),
      .dma_write_ctrl_rsci_bdwt(dma_write_ctrl_rsci_bdwt),
      .dma_write_ctrl_rsci_bcwt(dma_write_ctrl_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1 (
  clk, rst, plm_outputs_rsci_q_d, plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      core_wen, core_wten, plm_outputs_rsci_oswt_unreg, plm_outputs_rsci_bawt, plm_outputs_rsci_iswt0,
      plm_outputs_rsci_q_d_mxwt, plm_outputs_rsci_iswt0_pff
);
  input clk;
  input rst;
  input [31:0] plm_outputs_rsci_q_d;
  output plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input core_wen;
  input core_wten;
  input plm_outputs_rsci_oswt_unreg;
  output plm_outputs_rsci_bawt;
  input plm_outputs_rsci_iswt0;
  output [31:0] plm_outputs_rsci_q_d_mxwt;
  input plm_outputs_rsci_iswt0_pff;


  // Interconnect Declarations
  wire plm_outputs_rsci_biwt;
  wire plm_outputs_rsci_bdwt;
  wire plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl
      store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_ctrl_inst (
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsci_oswt_unreg(plm_outputs_rsci_oswt_unreg),
      .plm_outputs_rsci_iswt0(plm_outputs_rsci_iswt0),
      .plm_outputs_rsci_biwt(plm_outputs_rsci_biwt),
      .plm_outputs_rsci_bdwt(plm_outputs_rsci_bdwt),
      .plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct(plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct),
      .plm_outputs_rsci_iswt0_pff(plm_outputs_rsci_iswt0_pff)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp
      store_core_plm_outputs_rsci_1_plm_outputs_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsci_q_d(plm_outputs_rsci_q_d),
      .plm_outputs_rsci_bawt(plm_outputs_rsci_bawt),
      .plm_outputs_rsci_q_d_mxwt(plm_outputs_rsci_q_d_mxwt),
      .plm_outputs_rsci_biwt(plm_outputs_rsci_biwt),
      .plm_outputs_rsci_bdwt(plm_outputs_rsci_bdwt)
    );
  assign plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, core_wen, conf_info_rsci_oswt_unreg,
      conf_info_rsci_bawt, conf_info_rsci_iswt0, conf_info_rsci_wen_comp, conf_info_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input core_wen;
  input conf_info_rsci_oswt_unreg;
  output conf_info_rsci_bawt;
  input conf_info_rsci_iswt0;
  output conf_info_rsci_wen_comp;
  output [63:0] conf_info_rsci_idat_mxwt;


  // Interconnect Declarations
  wire conf_info_rsci_biwt;
  wire conf_info_rsci_bdwt;
  wire conf_info_rsci_bcwt;
  wire conf_info_rsci_irdy_core_sct;
  wire conf_info_rsci_ivld;
  wire [255:0] conf_info_rsci_idat;
  wire [63:0] conf_info_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_ccs_in_wait_v1 #(.rscid(32'sd23),
  .width(32'sd256)) conf_info_rsci (
      .rdy(conf_info_rsc_rdy),
      .vld(conf_info_rsc_vld),
      .dat(conf_info_rsc_dat),
      .irdy(conf_info_rsci_irdy_core_sct),
      .ivld(conf_info_rsci_ivld),
      .idat(conf_info_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_ctrl store_core_conf_info_rsci_conf_info_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_iswt0(conf_info_rsci_iswt0),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_irdy_core_sct(conf_info_rsci_irdy_core_sct),
      .conf_info_rsci_ivld(conf_info_rsci_ivld)
    );
  esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci_conf_info_wait_dp store_core_conf_info_rsci_conf_info_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsci_oswt_unreg(conf_info_rsci_oswt_unreg),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt_pconst),
      .conf_info_rsci_biwt(conf_info_rsci_biwt),
      .conf_info_rsci_bdwt(conf_info_rsci_bdwt),
      .conf_info_rsci_bcwt(conf_info_rsci_bcwt),
      .conf_info_rsci_idat(conf_info_rsci_idat)
    );
  assign conf_info_rsci_idat_mxwt = conf_info_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core (
  clk, rst, acc_done_rsc_vld, config_done_cns_rdy, config_done_cns_vld, load_done_cns_rdy,
      load_done_cns_vld, compute_done_cns_rdy, compute_done_cns_vld, store_done_cns_rdy,
      store_done_cns_vld
);
  input clk;
  input rst;
  output acc_done_rsc_vld;
  output config_done_cns_rdy;
  input config_done_cns_vld;
  output load_done_cns_rdy;
  input load_done_cns_vld;
  output compute_done_cns_rdy;
  input compute_done_cns_vld;
  output store_done_cns_rdy;
  input store_done_cns_vld;


  // Interconnect Declarations
  wire core_wen;
  wire acc_done_rsci_bawt;
  wire core_wten;
  wire config_done_cnsi_bawt;
  wire config_done_cnsi_wen_comp;
  wire load_done_cnsi_bawt;
  wire load_done_cnsi_wen_comp;
  reg load_done_cnsi_irdy_core_psct;
  wire compute_done_cnsi_bawt;
  wire compute_done_cnsi_wen_comp;
  wire store_done_cnsi_bawt;
  wire store_done_cnsi_wen_comp;
  wire [1:0] fsm_output;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_5;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_21;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_56_cse;
  reg main_stage_v_4;
  reg reg_store_done_cnsi_irdy_core_psct_cse;
  reg reg_compute_done_cnsi_irdy_core_psct_cse;
  reg reg_store_done_cnsi_oswt_cse;
  reg reg_load_done_cnsi_iswt0_cse;
  wire or_20_cse;
  wire or_17_cse;
  wire or_15_cse;
  wire or_cse;
  wire main_stage_v_4_mx0c1;
  reg reg_config_done_cnsi_iswt0_cse;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_acc_done_rsci conv2d_cxx_catapult_core_core_acc_done_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .acc_done_rsc_vld(acc_done_rsc_vld),
      .core_wen(core_wen),
      .acc_done_rsci_oswt_unreg(and_dcpl_27),
      .acc_done_rsci_bawt(acc_done_rsci_bawt),
      .acc_done_rsci_iswt0(reg_store_done_cnsi_oswt_cse),
      .core_wten(core_wten)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_config_done_cnsi conv2d_cxx_catapult_core_core_config_done_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .config_done_cns_rdy(config_done_cns_rdy),
      .config_done_cns_vld(config_done_cns_vld),
      .core_wen(core_wen),
      .config_done_cnsi_oswt_unreg(and_56_cse),
      .config_done_cnsi_bawt(config_done_cnsi_bawt),
      .config_done_cnsi_iswt0(reg_config_done_cnsi_iswt0_cse),
      .config_done_cnsi_wen_comp(config_done_cnsi_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_load_done_cnsi conv2d_cxx_catapult_core_core_load_done_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .load_done_cns_rdy(load_done_cns_rdy),
      .load_done_cns_vld(load_done_cns_vld),
      .core_wen(core_wen),
      .load_done_cnsi_oswt_unreg(and_dcpl_19),
      .load_done_cnsi_bawt(load_done_cnsi_bawt),
      .load_done_cnsi_iswt0(reg_load_done_cnsi_iswt0_cse),
      .load_done_cnsi_wen_comp(load_done_cnsi_wen_comp),
      .load_done_cnsi_irdy_core_psct(load_done_cnsi_irdy_core_psct)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_compute_done_cnsi conv2d_cxx_catapult_core_core_compute_done_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_done_cns_rdy(compute_done_cns_rdy),
      .compute_done_cns_vld(compute_done_cns_vld),
      .core_wen(core_wen),
      .compute_done_cnsi_oswt_unreg(and_dcpl_14),
      .compute_done_cnsi_bawt(compute_done_cnsi_bawt),
      .compute_done_cnsi_iswt0(reg_compute_done_cnsi_irdy_core_psct_cse),
      .compute_done_cnsi_wen_comp(compute_done_cnsi_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_store_done_cnsi conv2d_cxx_catapult_core_core_store_done_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .store_done_cns_rdy(store_done_cns_rdy),
      .store_done_cns_vld(store_done_cns_vld),
      .core_wen(core_wen),
      .store_done_cnsi_oswt_unreg(and_dcpl_18),
      .store_done_cnsi_bawt(store_done_cnsi_bawt),
      .store_done_cnsi_iswt0(reg_store_done_cnsi_irdy_core_psct_cse),
      .store_done_cnsi_wen_comp(store_done_cnsi_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_staller conv2d_cxx_catapult_core_core_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .config_done_cnsi_wen_comp(config_done_cnsi_wen_comp),
      .load_done_cnsi_wen_comp(load_done_cnsi_wen_comp),
      .compute_done_cnsi_wen_comp(compute_done_cnsi_wen_comp),
      .store_done_cnsi_wen_comp(store_done_cnsi_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core_core_fsm conv2d_cxx_catapult_core_core_core_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_20_cse = load_done_cnsi_bawt | (~ reg_load_done_cnsi_iswt0_cse);
  assign or_17_cse = compute_done_cnsi_bawt | (~ reg_compute_done_cnsi_irdy_core_psct_cse);
  assign or_15_cse = store_done_cnsi_bawt | (~ reg_store_done_cnsi_irdy_core_psct_cse);
  assign or_cse = acc_done_rsci_bawt | (~ main_stage_v_4);
  assign and_dcpl_1 = or_cse & or_15_cse;
  assign and_dcpl_2 = and_dcpl_1 & or_17_cse;
  assign and_dcpl_5 = load_done_cnsi_bawt & reg_load_done_cnsi_iswt0_cse;
  assign and_dcpl_13 = compute_done_cnsi_bawt & reg_compute_done_cnsi_irdy_core_psct_cse;
  assign and_dcpl_14 = and_dcpl_1 & and_dcpl_13;
  assign and_dcpl_17 = or_cse & store_done_cnsi_bawt & (~(compute_done_cnsi_bawt
      & reg_compute_done_cnsi_irdy_core_psct_cse)) & reg_store_done_cnsi_irdy_core_psct_cse;
  assign and_dcpl_18 = or_cse & reg_store_done_cnsi_irdy_core_psct_cse & store_done_cnsi_bawt;
  assign and_dcpl_19 = and_dcpl_2 & and_dcpl_5;
  assign and_dcpl_21 = and_dcpl_1 & and_dcpl_13 & (~(load_done_cnsi_bawt & reg_load_done_cnsi_iswt0_cse));
  assign and_dcpl_26 = and_dcpl_2 & and_dcpl_5 & (~ config_done_cnsi_bawt);
  assign and_dcpl_27 = main_stage_v_4 & acc_done_rsci_bawt;
  assign and_56_cse = and_dcpl_2 & or_20_cse & config_done_cnsi_bawt & (fsm_output[1]);
  assign main_stage_v_4_mx0c1 = and_dcpl_27 & (~(store_done_cnsi_bawt & reg_store_done_cnsi_irdy_core_psct_cse));
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_config_done_cnsi_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((config_done_cnsi_bawt & or_20_cse & or_17_cse & or_15_cse
        & or_cse) | (fsm_output[0])) ) begin
      reg_config_done_cnsi_iswt0_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_store_done_cnsi_irdy_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_14 | and_dcpl_17) ) begin
      reg_store_done_cnsi_irdy_core_psct_cse <= ~ and_dcpl_17;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_store_done_cnsi_oswt_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_store_done_cnsi_oswt_cse <= and_dcpl_18;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_compute_done_cnsi_irdy_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_19 | and_dcpl_21) ) begin
      reg_compute_done_cnsi_irdy_core_psct_cse <= ~ and_dcpl_21;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      load_done_cnsi_irdy_core_psct <= 1'b0;
    end
    else if ( core_wen & (and_56_cse | (and_dcpl_2 & and_dcpl_5 & config_done_cnsi_bawt)
        | and_dcpl_26) ) begin
      load_done_cnsi_irdy_core_psct <= ~ and_dcpl_26;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_load_done_cnsi_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (and_56_cse | and_dcpl_26) ) begin
      reg_load_done_cnsi_iswt0_cse <= ~ and_dcpl_26;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_18 | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config_core
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_conf_load_rsc_dat,
      plm_conf_load_rsc_vld, plm_conf_load_rsc_rdy, plm_conf_compute_rsc_dat, plm_conf_compute_rsc_vld,
      plm_conf_compute_rsc_rdy, plm_conf_store_rsc_dat, plm_conf_store_rsc_vld, plm_conf_store_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [255:0] plm_conf_load_rsc_dat;
  output plm_conf_load_rsc_vld;
  input plm_conf_load_rsc_rdy;
  output [255:0] plm_conf_compute_rsc_dat;
  output plm_conf_compute_rsc_vld;
  input plm_conf_compute_rsc_rdy;
  output [255:0] plm_conf_store_rsc_dat;
  output plm_conf_store_rsc_vld;
  input plm_conf_store_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire core_wen;
  wire conf_info_rsci_bawt;
  wire conf_info_rsci_wen_comp;
  wire [255:0] conf_info_rsci_idat_mxwt;
  wire plm_conf_load_rsci_bawt;
  wire plm_conf_load_rsci_wen_comp;
  wire plm_conf_compute_rsci_bawt;
  wire plm_conf_compute_rsci_wen_comp;
  wire plm_conf_store_rsci_bawt;
  wire plm_conf_store_rsci_wen_comp;
  reg [255:0] plm_conf_store_rsci_idat;
  wire done_rsci_bawt;
  wire done_rsci_wen_comp;
  wire [1:0] fsm_output;
  wire and_dcpl_1;
  wire and_dcpl_9;
  wire or_dcpl_3;
  wire or_dcpl_5;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire or_dcpl_6;
  wire and_dcpl_17;
  wire and_dcpl_20;
  wire or_tmp_8;
  reg reg_done_rsci_ivld_core_psct_cse;
  reg reg_plm_conf_store_rsci_ivld_core_psct_cse;
  reg [255:0] reg_plm_conf_compute_rsci_idat_cse;
  wire or_cse;
  reg reg_conf_info_rsci_iswt0_cse;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_config_core_conf_info_rsci config_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(or_tmp_8),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_iswt0(reg_conf_info_rsci_iswt0_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_load_rsci config_core_plm_conf_load_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_conf_load_rsc_dat(plm_conf_load_rsc_dat),
      .plm_conf_load_rsc_vld(plm_conf_load_rsc_vld),
      .plm_conf_load_rsc_rdy(plm_conf_load_rsc_rdy),
      .core_wen(core_wen),
      .plm_conf_load_rsci_oswt_unreg(and_dcpl_15),
      .plm_conf_load_rsci_bawt(plm_conf_load_rsci_bawt),
      .plm_conf_load_rsci_iswt0(reg_plm_conf_store_rsci_ivld_core_psct_cse),
      .plm_conf_load_rsci_wen_comp(plm_conf_load_rsci_wen_comp),
      .plm_conf_load_rsci_idat(reg_plm_conf_compute_rsci_idat_cse)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_compute_rsci config_core_plm_conf_compute_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_conf_compute_rsc_dat(plm_conf_compute_rsc_dat),
      .plm_conf_compute_rsc_vld(plm_conf_compute_rsc_vld),
      .plm_conf_compute_rsc_rdy(plm_conf_compute_rsc_rdy),
      .core_wen(core_wen),
      .plm_conf_compute_rsci_oswt_unreg(and_dcpl_15),
      .plm_conf_compute_rsci_bawt(plm_conf_compute_rsci_bawt),
      .plm_conf_compute_rsci_iswt0(reg_plm_conf_store_rsci_ivld_core_psct_cse),
      .plm_conf_compute_rsci_wen_comp(plm_conf_compute_rsci_wen_comp),
      .plm_conf_compute_rsci_idat(reg_plm_conf_compute_rsci_idat_cse)
    );
  esp_acc_conv2d_cxx_catapult_config_core_plm_conf_store_rsci config_core_plm_conf_store_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_conf_store_rsc_dat(plm_conf_store_rsc_dat),
      .plm_conf_store_rsc_vld(plm_conf_store_rsc_vld),
      .plm_conf_store_rsc_rdy(plm_conf_store_rsc_rdy),
      .core_wen(core_wen),
      .plm_conf_store_rsci_oswt_unreg(and_dcpl_15),
      .plm_conf_store_rsci_bawt(plm_conf_store_rsci_bawt),
      .plm_conf_store_rsci_iswt0(reg_plm_conf_store_rsci_ivld_core_psct_cse),
      .plm_conf_store_rsci_wen_comp(plm_conf_store_rsci_wen_comp),
      .plm_conf_store_rsci_idat(plm_conf_store_rsci_idat)
    );
  esp_acc_conv2d_cxx_catapult_config_core_done_rsci config_core_done_rsci_inst (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(and_dcpl_16),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_iswt0(reg_done_rsci_ivld_core_psct_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_config_core_staller config_core_staller_inst (
      .core_wen(core_wen),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .plm_conf_load_rsci_wen_comp(plm_conf_load_rsci_wen_comp),
      .plm_conf_compute_rsci_wen_comp(plm_conf_compute_rsci_wen_comp),
      .plm_conf_store_rsci_wen_comp(plm_conf_store_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_config_core_core_fsm config_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_cse = done_rsci_bawt | (~ reg_done_rsci_ivld_core_psct_cse);
  assign and_dcpl_1 = plm_conf_load_rsci_bawt & plm_conf_compute_rsci_bawt;
  assign and_dcpl_9 = reg_done_rsci_ivld_core_psct_cse & (~ done_rsci_bawt);
  assign or_dcpl_3 = ~(plm_conf_load_rsci_bawt & plm_conf_compute_rsci_bawt);
  assign or_dcpl_5 = ((or_dcpl_3 | (~ plm_conf_store_rsci_bawt)) & reg_plm_conf_store_rsci_ivld_core_psct_cse)
      | and_dcpl_9 | (~ conf_info_rsci_bawt);
  assign and_dcpl_15 = or_cse & plm_conf_load_rsci_bawt & plm_conf_compute_rsci_bawt
      & plm_conf_store_rsci_bawt & reg_plm_conf_store_rsci_ivld_core_psct_cse;
  assign and_dcpl_16 = reg_done_rsci_ivld_core_psct_cse & done_rsci_bawt;
  assign or_dcpl_6 = ~(plm_conf_store_rsci_bawt & reg_plm_conf_store_rsci_ivld_core_psct_cse);
  assign and_dcpl_17 = (or_dcpl_3 | or_dcpl_6) & and_dcpl_16;
  assign and_dcpl_20 = or_cse & and_dcpl_1 & plm_conf_store_rsci_bawt & reg_plm_conf_store_rsci_ivld_core_psct_cse
      & (~ conf_info_rsci_bawt);
  assign or_tmp_8 = (~((~(and_dcpl_1 & plm_conf_store_rsci_bawt)) & reg_plm_conf_store_rsci_ivld_core_psct_cse))
      & or_cse & conf_info_rsci_bawt & (fsm_output[1]);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((conf_info_rsci_bawt & (plm_conf_load_rsci_bawt | (~ reg_plm_conf_store_rsci_ivld_core_psct_cse))
        & (plm_conf_compute_rsci_bawt | (~ reg_plm_conf_store_rsci_ivld_core_psct_cse))
        & (plm_conf_store_rsci_bawt | (~ reg_plm_conf_store_rsci_ivld_core_psct_cse))
        & or_cse) | (fsm_output[0])) ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_done_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_15 | and_dcpl_17) ) begin
      reg_done_rsci_ivld_core_psct_cse <= ~ and_dcpl_17;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_conf_store_rsci_idat <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_5 | ((and_dcpl_9 | or_dcpl_3 | or_dcpl_6 | (~
        conf_info_rsci_bawt)) & (fsm_output[0])))) ) begin
      plm_conf_store_rsci_idat <= conf_info_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_conf_store_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (or_tmp_8 | and_dcpl_20) ) begin
      reg_plm_conf_store_rsci_ivld_core_psct_cse <= ~ and_dcpl_20;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_conf_compute_rsci_idat_cse <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~(or_dcpl_5 | (fsm_output[0]))) ) begin
      reg_plm_conf_compute_rsci_idat_cse <= conf_info_rsci_idat_mxwt;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load_core
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_inputs_rsc_req_vz,
      plm_inputs_rsc_rls_lz, plm_filters_rsc_req_vz, plm_filters_rsc_rls_lz, dma_read_ctrl_rsc_dat,
      dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld,
      dma_read_chnl_rsc_rdy, done_rsc_rdy, done_rsc_vld, plm_inputs_rsci_d_d, plm_inputs_rsci_wadr_d,
      plm_filters_rsci_d_d, plm_filters_rsci_wadr_d, plm_inputs_rsci_we_d_pff, plm_filters_rsci_we_d_pff
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input plm_inputs_rsc_req_vz;
  output plm_inputs_rsc_rls_lz;
  input plm_filters_rsc_req_vz;
  output plm_filters_rsc_rls_lz;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;
  output [31:0] plm_inputs_rsci_d_d;
  output [13:0] plm_inputs_rsci_wadr_d;
  output [31:0] plm_filters_rsci_d_d;
  output [15:0] plm_filters_rsci_wadr_d;
  output plm_inputs_rsci_we_d_pff;
  output plm_filters_rsci_we_d_pff;


  // Interconnect Declarations
  wire core_wen;
  wire conf_info_rsci_bawt;
  wire core_wten;
  wire conf_info_rsci_wen_comp;
  wire [63:0] conf_info_rsci_idat_mxwt;
  wire plm_inputs_rsci_bawt;
  wire plm_filters_rsci_bawt;
  wire dma_read_ctrl_rsci_bawt;
  wire dma_read_ctrl_rsci_irdy_mxwt;
  wire dma_read_chnl_rsci_bawt;
  wire dma_read_chnl_rsci_wen_comp;
  wire [31:0] dma_read_chnl_rsci_idat_mxwt;
  wire done_rsci_bawt;
  wire done_rsci_wen_comp;
  wire plm_inputs_rsc_rls_obj_bawt;
  wire plm_filters_rsc_rls_obj_bawt;
  wire plm_inputs_rsc_req_obj_bawt;
  wire plm_inputs_rsc_req_obj_wen_comp;
  wire plm_filters_rsc_req_obj_bawt;
  wire plm_filters_rsc_req_obj_wen_comp;
  reg [15:0] dma_read_ctrl_rsci_idat_47_32;
  reg [15:0] dma_read_ctrl_rsci_idat_15_0;
  wire [1:0] fsm_output;
  wire LOAD_LOOP_LOAD_LOOP_if_and_tmp;
  wire LOAD_BATCH_LOOP_if_1_equal_tmp;
  wire [8:0] operator_8_false_4_acc_tmp;
  wire [9:0] nl_operator_8_false_4_acc_tmp;
  wire [5:0] PADDING_LOOP_acc_tmp;
  wire [6:0] nl_PADDING_LOOP_acc_tmp;
  wire PADDING_LOOP_if_equal_tmp;
  wire [8:0] operator_8_false_3_acc_tmp;
  wire [9:0] nl_operator_8_false_3_acc_tmp;
  wire PADDING_LOOP_for_if_equal_tmp;
  wire [8:0] operator_8_false_2_acc_tmp;
  wire [9:0] nl_operator_8_false_2_acc_tmp;
  wire PADDING_LOOP_for_for_if_1_equal_tmp;
  wire [8:0] operator_8_false_1_acc_tmp;
  wire [9:0] nl_operator_8_false_1_acc_tmp;
  wire and_7_tmp;
  wire and_5_tmp;
  wire and_3_tmp;
  wire or_tmp_3;
  wire or_tmp_10;
  wire or_tmp_18;
  wire or_tmp_64;
  wire mux_tmp_65;
  wire or_tmp_86;
  wire and_dcpl_1;
  wire or_tmp_92;
  wire not_tmp_61;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire or_tmp_109;
  wire mux_tmp_76;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_19;
  wire and_dcpl_22;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire or_dcpl_18;
  wire or_dcpl_19;
  wire mux_tmp_85;
  wire not_tmp_85;
  wire or_dcpl_23;
  wire or_dcpl_25;
  wire mux_tmp_95;
  wire and_dcpl_54;
  wire or_dcpl_39;
  wire or_tmp_137;
  wire or_tmp_152;
  wire PADDING_LOOP_mux_11_cse;
  wire and_165_cse;
  wire [4:0] LOAD_BATCH_LOOP_b_4_0_sva_2;
  wire [5:0] nl_LOAD_BATCH_LOOP_b_4_0_sva_2;
  wire exit_PADDING_LOOP_lpi_1_dfm_2_mx1;
  wire PADDING_LOOP_equal_tmp_1_mx0w0;
  wire [15:0] LOAD_LOOP_i_lpi_1_mx0;
  wire [32:0] operator_32_false_acc_psp_sva_1;
  wire [33:0] nl_operator_32_false_acc_psp_sva_1;
  wire exit_PADDING_LOOP_for_lpi_1_dfm_4;
  wire exit_PADDING_LOOP_sva_2;
  wire exit_PADDING_LOOP_for_for_lpi_1_dfm_1;
  wire exit_PADDING_LOOP_for_sva_5;
  wire lfst_exit_PADDING_LOOP_lpi_1_dfm_1_mx0w0;
  wire lfst_exit_PADDING_LOOP_lpi_1_dfm_0_mx0w0;
  wire exitL_exit_PADDING_LOOP_lpi_1_mx0;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_3;
  reg exitL_exit_LOAD_BATCH_LOOP_sva;
  wire lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1_mx0w0;
  wire lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0_mx0w0;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0;
  reg PADDING_LOOP_equal_tmp_1_1;
  wire PADDING_LOOP_and_2_ssc_1;
  reg PADDING_LOOP_or_tmp_1;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_3;
  reg main_stage_v_3;
  reg lfst_exit_PADDING_LOOP_for_1_lpi_1;
  wire PADDING_LOOP_or_tmp_mx0w0;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0;
  reg exitL_exit_PADDING_LOOP_lpi_1;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_2_1_0;
  reg exit_LOAD_LOOP_sva_1;
  reg PADDING_LOOP_equal_tmp_1;
  reg LOAD_BATCH_LOOP_asn_itm;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1;
  reg exit_LOAD_CTRL_LOOP_sva_st_1;
  reg exit_PADDING_LOOP_lpi_1_dfm_2_st_1;
  reg lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0;
  reg exit_PADDING_LOOP_lpi_1_dfm_2_st_2;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_2;
  reg PADDING_LOOP_for_for_land_2_lpi_1_dfm_st_1;
  wire exit_LOAD_BATCH_LOOP_sva_2_mx0w0;
  reg exit_LOAD_BATCH_LOOP_sva_2;
  wire exit_PADDING_LOOP_lpi_1_dfm_mx0w0;
  reg exit_PADDING_LOOP_lpi_1_dfm;
  wire exit_PADDING_LOOP_for_lpi_1_dfm_1_mx0w0;
  reg exit_PADDING_LOOP_for_lpi_1_dfm_1;
  wire exit_LOAD_LOOP_lpi_1_dfm_mx1w0;
  wire PADDING_LOOP_equal_tmp_mx1w0;
  wire exitL_exit_PADDING_LOOP_lpi_1_dfm_1;
  reg reg_conf_info_rsci_iswt0_cse;
  reg reg_plm_filters_rsc_req_obj_iswt0_cse;
  reg reg_plm_filters_rsc_rls_obj_ld_core_psct_cse;
  reg reg_done_rsci_ivld_core_psct_cse;
  reg reg_dma_read_chnl_rsci_irdy_core_psct_cse;
  reg reg_dma_read_ctrl_rsci_ivld_core_psct_cse;
  reg reg_plm_filters_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse;
  reg reg_plm_inputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse;
  wire PADDING_LOOP_and_cse;
  wire and_193_cse;
  wire LOAD_BATCH_LOOP_and_cse;
  wire or_38_cse;
  wire PADDING_LOOP_and_17_cse;
  wire or_62_cse;
  wire or_42_cse;
  wire or_73_cse;
  wire or_162_cse;
  wire PADDING_LOOP_nor_cse;
  wire and_115_cse;
  wire mux_70_cse;
  wire and_197_cse;
  wire nor_24_cse;
  reg [31:0] plm_inputs_rsci_d_d_reg;
  wire [31:0] PADDING_LOOP_for_for_mux_rmff;
  reg [13:0] plm_inputs_rsci_wadr_d_reg;
  wire [13:0] PADDING_LOOP_for_for_index_in_mux_rmff;
  wire plm_inputs_rsci_we_d_iff;
  wire and_60_rmff;
  reg [31:0] plm_filters_rsci_d_d_reg;
  wire [31:0] LOAD_LOOP_data_ac_mux_rmff;
  reg [15:0] plm_filters_rsci_wadr_d_reg;
  wire [15:0] LOAD_LOOP_i_mux_rmff;
  wire plm_filters_rsci_we_d_iff;
  wire and_58_rmff;
  wire and_42_rmff;
  wire and_dcpl_58;
  wire PADDING_LOOP_for_for_and_3_psp_mx1;
  wire PADDING_LOOP_and_8_m1c_1;
  wire PADDING_LOOP_for_for_and_3_psp_mx1w0;
  reg [4:0] PADDING_LOOP_for_row_4_0_lpi_1;
  wire [4:0] PADDING_LOOP_for_row_4_0_sva_2;
  wire [5:0] nl_PADDING_LOOP_for_row_4_0_sva_2;
  wire or_296_tmp;
  wire PADDING_LOOP_and_3_tmp;
  wire and_219_cse;
  wire [15:0] z_out;
  wire [23:0] nl_z_out;
  wire [15:0] z_out_1;
  wire [23:0] nl_z_out_1;
  wire [15:0] z_out_2;
  wire [23:0] nl_z_out_2;
  reg [15:0] LOAD_LOOP_i_lpi_1;
  reg [4:0] PADDING_LOOP_for_for_col_4_0_lpi_1;
  reg [7:0] pad_lpi_1_dfm;
  reg [15:0] ac_int_cctor_8_lpi_1_dfm;
  reg [6:0] n_w_in_acc_psp_lpi_1_dfm;
  wire [7:0] nl_n_w_in_acc_psp_lpi_1_dfm;
  reg [6:0] n_h_in_acc_psp_lpi_1_dfm;
  wire [7:0] nl_n_h_in_acc_psp_lpi_1_dfm;
  reg [15:0] mul_4_cse_lpi_1_dfm;
  reg [15:0] LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm;
  reg PADDING_LOOP_for_and_psp;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg exit_LOAD_CTRL_LOOP_sva_st;
  reg PADDING_LOOP_for_for_land_2_lpi_1_dfm_st;
  reg [15:0] LOAD_LOOP_i_sva_1_1;
  reg PADDING_LOOP_for_for_land_2_lpi_1_dfm_1;
  reg [13:0] PADDING_LOOP_for_for_index_in_acc_itm_1;
  wire [14:0] nl_PADDING_LOOP_for_for_index_in_acc_itm_1;
  reg [3:0] LOAD_BATCH_LOOP_b_4_0_lpi_1_3_0;
  reg [4:0] PADDING_LOOP_chan_5_0_lpi_1_4_0;
  reg [7:0] conf_info_crt_lpi_1_dfm_231_224;
  reg conf_info_crt_lpi_1_dfm_192;
  reg conf_info_crt_lpi_1_dfm_160;
  reg [7:0] conf_info_crt_lpi_1_dfm_135_128;
  reg [7:0] conf_info_crt_lpi_1_dfm_71_64;
  reg PADDING_LOOP_for_for_and_3_psp;
  wire [15:0] LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm_mx0w0;
  wire [19:0] nl_LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm_mx0w0;
  wire dma_read_ctrl_rsci_idat_15_0_mx0c1;
  wire dma_read_ctrl_rsci_idat_47_32_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire [15:0] ac_int_cctor_8_lpi_1_dfm_mx0;
  wire exit_PADDING_LOOP_lpi_1_dfm_2_mx1w0;
  wire main_stage_v_1_mx0c1;
  wire [15:0] LOAD_LOOP_i_sva_1_mx0w0;
  wire [16:0] nl_LOAD_LOOP_i_sva_1_mx0w0;
  wire exit_PADDING_LOOP_lpi_1_dfm_2_st_1_mx0c1;
  wire PADDING_LOOP_for_for_land_2_lpi_1_dfm_mx0w0;
  wire exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_mx0w0;
  wire PADDING_LOOP_for_and_psp_mx1w0;
  wire [3:0] LOAD_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1;
  wire [4:0] PADDING_LOOP_for_for_col_4_0_lpi_1_dfm_3;
  wire [4:0] PADDING_LOOP_for_for_col_4_0_sva_2;
  wire [5:0] nl_PADDING_LOOP_for_for_col_4_0_sva_2;
  wire [15:0] ac_int_cctor_8_sva_1;
  wire [16:0] nl_ac_int_cctor_8_sva_1;
  wire [15:0] mul_4_cse_sva_1;
  wire [7:0] pad_sva_1;
  wire signed [16:0] nl_pad_sva_1;
  wire or_10_cse_1;
  wire or_11_cse_1;
  wire or_12_cse_1;
  wire or_13_cse_1;
  wire or_4_cse_1;
  wire or_5_cse_1;
  wire or_6_cse_1;
  wire or_cse_1;
  wire nand_21_cse_1;
  wire PADDING_LOOP_or_cse_1;
  wire nand_5_cse_1;
  wire nand_9_cse_1;
  wire [16:0] pad_acc_psp_sva_1;
  wire [17:0] nl_pad_acc_psp_sva_1;
  wire PADDING_LOOP_for_for_aelse_acc_itm_8;
  wire PADDING_LOOP_and_7_rgt;
  wire PADDING_LOOP_and_11_rgt;
  wire and_73_rgt;
  wire and_223_cse;
  wire and_234_cse;
  wire LOAD_LOOP_and_cse;
  wire LOAD_LOOP_i_and_cse;
  wire PADDING_LOOP_and_31_cse;
  reg reg_exit_PADDING_LOOP_lpi_1_dfm_2_cse;
  wire PADDING_LOOP_for_for_aelse_2_acc_itm_9_1;
  wire PADDING_LOOP_for_for_aelse_1_acc_itm_9_1;
  wire operator_8_false_2_acc_itm_4_1;
  wire operator_8_false_3_acc_itm_4_1;
  wire PADDING_LOOP_for_for_if_acc_itm_8;

  wire[0:0] or_61_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] and_53_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] nand_48_nl;
  wire[0:0] nor_13_nl;
  wire[31:0] PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] PADDING_LOOP_for_row_PADDING_LOOP_for_row_PADDING_LOOP_for_row_mux_nl;
  wire[0:0] PADDING_LOOP_and_9_nl;
  wire[0:0] and_217_nl;
  wire[0:0] PADDING_LOOP_for_mux_4_nl;
  wire[0:0] LOAD_LOOP_LOAD_LOOP_and_2_nl;
  wire[12:0] PADDING_LOOP_for_for_index_in_acc_2_nl;
  wire[13:0] nl_PADDING_LOOP_for_for_index_in_acc_2_nl;
  wire[0:0] nor_47_nl;
  wire[0:0] and_221_nl;
  wire[0:0] PADDING_LOOP_mux_7_nl;
  wire[0:0] or_201_nl;
  wire[0:0] PADDING_LOOP_PADDING_LOOP_nor_nl;
  wire[6:0] operator_16_false_acc_nl;
  wire[7:0] nl_operator_16_false_acc_nl;
  wire[0:0] PADDING_LOOP_mux_10_nl;
  wire[0:0] PADDING_LOOP_mux_13_nl;
  wire[0:0] LOAD_BATCH_LOOP_mux_8_nl;
  wire[31:0] LOAD_LOOP_mul_nl;
  wire[23:0] LOAD_LOOP_mul_1_nl;
  wire[0:0] LOAD_BATCH_LOOP_not_17_nl;
  wire[9:0] PADDING_LOOP_for_for_aelse_2_acc_nl;
  wire[10:0] nl_PADDING_LOOP_for_for_aelse_2_acc_nl;
  wire[8:0] PADDING_LOOP_for_for_aelse_2_acc_1_nl;
  wire[9:0] nl_PADDING_LOOP_for_for_aelse_2_acc_1_nl;
  wire[9:0] PADDING_LOOP_for_for_aelse_1_acc_nl;
  wire[10:0] nl_PADDING_LOOP_for_for_aelse_1_acc_nl;
  wire[8:0] PADDING_LOOP_for_for_aelse_1_acc_1_nl;
  wire[9:0] nl_PADDING_LOOP_for_for_aelse_1_acc_1_nl;
  wire[8:0] PADDING_LOOP_for_for_aelse_acc_nl;
  wire[9:0] nl_PADDING_LOOP_for_for_aelse_acc_nl;
  wire[4:0] operator_8_false_2_acc_nl;
  wire[5:0] nl_operator_8_false_2_acc_nl;
  wire[4:0] operator_8_false_3_acc_nl;
  wire[5:0] nl_operator_8_false_3_acc_nl;
  wire[0:0] PADDING_LOOP_for_mux_1_nl;
  wire[8:0] PADDING_LOOP_for_for_if_acc_nl;
  wire[9:0] nl_PADDING_LOOP_for_for_if_acc_nl;
  wire[7:0] operator_43_true_operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_operator_43_true_acc_nl;
  wire[0:0] operator_43_true_and_nl;
  wire[8:0] pad_acc_2_nl;
  wire[9:0] nl_pad_acc_2_nl;
  wire[16:0] pad_mul_nl;
  wire signed [17:0] nl_pad_mul_nl;
  wire[8:0] operator_8_false_acc_nl;
  wire[9:0] nl_operator_8_false_acc_nl;
  wire[0:0] or_115_nl;
  wire[0:0] or_50_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] nand_67_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] or_118_nl;
  wire[0:0] or_116_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] or_126_nl;
  wire[0:0] nor_40_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] or_196_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] or_205_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] nor_18_nl;
  wire[0:0] and_194_nl;
  wire[7:0] PADDING_LOOP_for_for_index_in_mux_8_nl;
  wire[15:0] PADDING_LOOP_for_for_index_in_mux_9_nl;
  wire[7:0] PADDING_LOOP_for_for_index_in_mux_10_nl;
  wire[15:0] PADDING_LOOP_for_for_index_in_mux_11_nl;
  wire[15:0] mul_6_nl;
  wire[7:0] PADDING_LOOP_for_for_index_in_mux_12_nl;
  wire[15:0] PADDING_LOOP_for_for_index_in_mux_13_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_load_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg;
  assign nl_load_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg = and_dcpl_1
      & (fsm_output[1]);
  wire [0:0] nl_load_core_plm_inputs_rsci_1_inst_plm_inputs_rsci_oswt_unreg;
  assign nl_load_core_plm_inputs_rsci_1_inst_plm_inputs_rsci_oswt_unreg = and_dcpl_22
      & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0;
  wire [0:0] nl_load_core_plm_filters_rsci_1_inst_plm_filters_rsci_oswt_unreg;
  assign nl_load_core_plm_filters_rsci_1_inst_plm_filters_rsci_oswt_unreg = and_dcpl_22
      & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0);
  wire [66:0] nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat;
  assign nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat = {19'b0110000000000000000
      , dma_read_ctrl_rsci_idat_47_32 , 16'b0000000000000000 , dma_read_ctrl_rsci_idat_15_0};
  wire [0:0] nl_load_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg;
  assign nl_load_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg = or_dcpl_18
      & and_dcpl_30;
  esp_acc_conv2d_cxx_catapult_load_core_conf_info_rsci load_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(nl_load_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg[0:0]),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_iswt0(reg_conf_info_rsci_iswt0_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsci_1 load_core_plm_inputs_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsci_oswt_unreg(nl_load_core_plm_inputs_rsci_1_inst_plm_inputs_rsci_oswt_unreg[0:0]),
      .plm_inputs_rsci_bawt(plm_inputs_rsci_bawt),
      .plm_inputs_rsci_iswt0(reg_plm_inputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse),
      .plm_inputs_rsci_we_d_pff(plm_inputs_rsci_we_d_iff),
      .plm_inputs_rsci_iswt0_pff(and_60_rmff)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsci_1 load_core_plm_filters_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsci_oswt_unreg(nl_load_core_plm_filters_rsci_1_inst_plm_filters_rsci_oswt_unreg[0:0]),
      .plm_filters_rsci_bawt(plm_filters_rsci_bawt),
      .plm_filters_rsci_iswt0(reg_plm_filters_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse),
      .plm_filters_rsci_we_d_pff(plm_filters_rsci_we_d_iff),
      .plm_filters_rsci_iswt0_pff(and_58_rmff)
    );
  esp_acc_conv2d_cxx_catapult_load_core_dma_read_ctrl_rsci load_core_dma_read_ctrl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .dma_read_ctrl_rsci_oswt_unreg(or_tmp_152),
      .dma_read_ctrl_rsci_bawt(dma_read_ctrl_rsci_bawt),
      .dma_read_ctrl_rsci_iswt0(reg_dma_read_ctrl_rsci_ivld_core_psct_cse),
      .dma_read_ctrl_rsci_irdy_mxwt(dma_read_ctrl_rsci_irdy_mxwt),
      .dma_read_ctrl_rsci_idat(nl_load_core_dma_read_ctrl_rsci_inst_dma_read_ctrl_rsci_idat[66:0])
    );
  esp_acc_conv2d_cxx_catapult_load_core_dma_read_chnl_rsci load_core_dma_read_chnl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .core_wen(core_wen),
      .dma_read_chnl_rsci_oswt_unreg(nl_load_core_dma_read_chnl_rsci_inst_dma_read_chnl_rsci_oswt_unreg[0:0]),
      .dma_read_chnl_rsci_bawt(dma_read_chnl_rsci_bawt),
      .dma_read_chnl_rsci_iswt0(reg_dma_read_chnl_rsci_irdy_core_psct_cse),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .dma_read_chnl_rsci_idat_mxwt(dma_read_chnl_rsci_idat_mxwt)
    );
  esp_acc_conv2d_cxx_catapult_load_core_done_rsci load_core_done_rsci_inst (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(and_dcpl_26),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_iswt0(reg_done_rsci_ivld_core_psct_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_rls_obj load_core_plm_inputs_rsc_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_rls_lz(plm_inputs_rsc_rls_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsc_rls_obj_oswt_unreg(and_42_rmff),
      .plm_inputs_rsc_rls_obj_bawt(plm_inputs_rsc_rls_obj_bawt),
      .plm_inputs_rsc_rls_obj_iswt0(reg_plm_filters_rsc_rls_obj_ld_core_psct_cse)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_rls_obj load_core_plm_filters_rsc_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_rls_lz(plm_filters_rsc_rls_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsc_rls_obj_oswt_unreg(and_42_rmff),
      .plm_filters_rsc_rls_obj_bawt(plm_filters_rsc_rls_obj_bawt),
      .plm_filters_rsc_rls_obj_iswt0(reg_plm_filters_rsc_rls_obj_ld_core_psct_cse)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_inputs_rsc_req_obj load_core_plm_inputs_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_req_vz(plm_inputs_rsc_req_vz),
      .core_wen(core_wen),
      .plm_inputs_rsc_req_obj_oswt_unreg(and_dcpl_15),
      .plm_inputs_rsc_req_obj_bawt(plm_inputs_rsc_req_obj_bawt),
      .plm_inputs_rsc_req_obj_iswt0(reg_plm_filters_rsc_req_obj_iswt0_cse),
      .plm_inputs_rsc_req_obj_wen_comp(plm_inputs_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_load_core_plm_filters_rsc_req_obj load_core_plm_filters_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_req_vz(plm_filters_rsc_req_vz),
      .core_wen(core_wen),
      .plm_filters_rsc_req_obj_oswt_unreg(and_dcpl_15),
      .plm_filters_rsc_req_obj_bawt(plm_filters_rsc_req_obj_bawt),
      .plm_filters_rsc_req_obj_iswt0(reg_plm_filters_rsc_req_obj_iswt0_cse),
      .plm_filters_rsc_req_obj_wen_comp(plm_filters_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_load_core_staller load_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .dma_read_chnl_rsci_wen_comp(dma_read_chnl_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .plm_inputs_rsc_req_obj_wen_comp(plm_inputs_rsc_req_obj_wen_comp),
      .plm_filters_rsc_req_obj_wen_comp(plm_filters_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_load_core_core_fsm load_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_61_nl = PADDING_LOOP_or_tmp_1 | (~ PADDING_LOOP_mux_11_cse);
  assign mux_70_cse = MUX_s_1_2_2(or_62_cse, or_61_nl, and_5_tmp);
  assign and_197_cse = ((~ PADDING_LOOP_for_for_if_1_equal_tmp) | (operator_8_false_1_acc_tmp[8:5]!=4'b0000))
      & operator_8_false_3_acc_itm_4_1;
  assign LOAD_BATCH_LOOP_and_cse = core_wen & (~((~ and_7_tmp) | (fsm_output[0])));
  assign and_42_rmff = and_dcpl_22 & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0 & exit_PADDING_LOOP_lpi_1_dfm_2_st_2;
  assign and_58_rmff = (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0) & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1
      & and_5_tmp;
  assign and_60_rmff = and_dcpl_19 & and_5_tmp;
  assign LOAD_LOOP_i_mux_rmff = MUX_v_16_2_2(LOAD_LOOP_i_lpi_1, plm_filters_rsci_wadr_d_reg,
      or_dcpl_23);
  assign LOAD_LOOP_data_ac_mux_rmff = MUX_v_32_2_2(dma_read_chnl_rsci_idat_mxwt,
      plm_filters_rsci_d_d_reg, or_dcpl_23);
  assign PADDING_LOOP_for_for_index_in_mux_rmff = MUX_v_14_2_2(PADDING_LOOP_for_for_index_in_acc_itm_1,
      plm_inputs_rsci_wadr_d_reg, or_dcpl_25);
  assign PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      dma_read_chnl_rsci_idat_mxwt, PADDING_LOOP_for_for_land_2_lpi_1_dfm_1);
  assign PADDING_LOOP_for_for_mux_rmff = MUX_v_32_2_2(PADDING_LOOP_for_for_PADDING_LOOP_for_for_and_nl,
      plm_inputs_rsci_d_d_reg, or_dcpl_25);
  assign and_115_cse = and_7_tmp & (fsm_output[1]);
  assign PADDING_LOOP_and_cse = core_wen & (~((~ and_5_tmp) | (fsm_output[0])));
  assign or_38_cse = (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1) | lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0
      | exitL_exit_PADDING_LOOP_lpi_1;
  assign or_42_cse = (~ PADDING_LOOP_equal_tmp_1_1) | lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0;
  assign and_234_cse = core_wen & exitL_exit_LOAD_BATCH_LOOP_sva;
  assign PADDING_LOOP_and_17_cse = core_wen & (~ (fsm_output[0]));
  assign PADDING_LOOP_and_31_cse = PADDING_LOOP_and_17_cse & (~(mux_70_cse | or_dcpl_19));
  assign and_193_cse = ((~ PADDING_LOOP_for_if_equal_tmp) | (operator_8_false_2_acc_tmp[8:5]!=4'b0000))
      & operator_8_false_2_acc_itm_4_1;
  assign PADDING_LOOP_for_mux_4_nl = MUX_s_1_2_2(PADDING_LOOP_for_and_psp_mx1w0,
      PADDING_LOOP_for_and_psp, or_dcpl_39);
  assign PADDING_LOOP_and_7_rgt = PADDING_LOOP_for_mux_4_nl & PADDING_LOOP_equal_tmp_1_mx0w0
      & and_7_tmp;
  assign PADDING_LOOP_and_11_rgt = exit_PADDING_LOOP_for_for_lpi_1_dfm_1 & PADDING_LOOP_equal_tmp_1_mx0w0
      & and_7_tmp;
  assign and_73_rgt = or_tmp_86 & and_7_tmp;
  assign LOAD_LOOP_i_and_cse = core_wen & and_7_tmp;
  assign LOAD_LOOP_and_cse = PADDING_LOOP_and_17_cse & and_7_tmp;
  assign nl_LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm_mx0w0 = ac_int_cctor_8_lpi_1_dfm_mx0
      * LOAD_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1;
  assign LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm_mx0w0 = nl_LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm_mx0w0[15:0];
  assign and_219_cse = (~ dma_read_ctrl_rsci_irdy_mxwt) & PADDING_LOOP_or_tmp_1;
  assign or_296_tmp = and_219_cse | PADDING_LOOP_equal_tmp_1_1 | (exit_LOAD_LOOP_sva_1
      & PADDING_LOOP_equal_tmp_1) | (~ and_5_tmp);
  assign PADDING_LOOP_and_3_tmp = (~ exit_LOAD_LOOP_sva_1) & PADDING_LOOP_equal_tmp_1
      & and_5_tmp;
  assign nor_47_nl = ~(PADDING_LOOP_and_3_tmp | or_296_tmp);
  assign and_221_nl = PADDING_LOOP_and_3_tmp & (~ or_296_tmp);
  assign LOAD_LOOP_i_lpi_1_mx0 = MUX1HOT_v_16_3_2((signext_16_1(~ dma_read_ctrl_rsci_irdy_mxwt)),
      LOAD_LOOP_i_sva_1_1, LOAD_LOOP_i_lpi_1, {nor_47_nl , and_221_nl , or_296_tmp});
  assign ac_int_cctor_8_lpi_1_dfm_mx0 = MUX_v_16_2_2(ac_int_cctor_8_lpi_1_dfm, ac_int_cctor_8_sva_1,
      exitL_exit_LOAD_BATCH_LOOP_sva);
  assign LOAD_BATCH_LOOP_if_1_equal_tmp = LOAD_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1 ==
      (operator_8_false_4_acc_tmp[3:0]);
  assign exit_LOAD_BATCH_LOOP_sva_2_mx0w0 = ~((~(LOAD_BATCH_LOOP_if_1_equal_tmp &
      (operator_8_false_4_acc_tmp[7:4]==4'b0000))) | (operator_8_false_4_acc_tmp[8]));
  assign or_201_nl = and_193_cse | and_197_cse;
  assign PADDING_LOOP_mux_7_nl = MUX_s_1_2_2(exit_PADDING_LOOP_lpi_1_dfm_mx0w0, exit_PADDING_LOOP_lpi_1_dfm,
      or_201_nl);
  assign exit_PADDING_LOOP_lpi_1_dfm_2_mx1w0 = PADDING_LOOP_mux_7_nl & exit_PADDING_LOOP_for_lpi_1_dfm_4;
  assign exit_PADDING_LOOP_lpi_1_dfm_2_mx1 = MUX_s_1_2_2(exit_PADDING_LOOP_lpi_1_dfm_2_mx1w0,
      reg_exit_PADDING_LOOP_lpi_1_dfm_2_cse, or_tmp_64);
  assign exit_PADDING_LOOP_lpi_1_dfm_mx0w0 = (PADDING_LOOP_acc_tmp[5]) | exit_PADDING_LOOP_sva_2;
  assign exit_PADDING_LOOP_for_lpi_1_dfm_1_mx0w0 = (~ operator_8_false_2_acc_itm_4_1)
      | exit_PADDING_LOOP_for_sva_5;
  assign PADDING_LOOP_PADDING_LOOP_nor_nl = ~(lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1_mx0w0
      | lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0_mx0w0);
  assign exitL_exit_PADDING_LOOP_lpi_1_mx0 = MUX_s_1_2_2(exitL_exit_PADDING_LOOP_lpi_1,
      PADDING_LOOP_PADDING_LOOP_nor_nl, and_5_tmp);
  assign PADDING_LOOP_nor_cse = ~(lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0 | (~ PADDING_LOOP_equal_tmp_1_1));
  assign lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1_mx0w0 = (~(PADDING_LOOP_nor_cse | and_219_cse))
      | PADDING_LOOP_and_2_ssc_1;
  assign PADDING_LOOP_mux_11_cse = MUX_s_1_2_2(lfst_exit_PADDING_LOOP_lpi_1_dfm_2_1_0,
      lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0, PADDING_LOOP_equal_tmp_1_1);
  assign lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0_mx0w0 = (PADDING_LOOP_mux_11_cse &
      (~ PADDING_LOOP_and_2_ssc_1)) | and_219_cse;
  assign PADDING_LOOP_or_tmp_mx0w0 = (lfst_exit_PADDING_LOOP_lpi_1_dfm_0_mx0w0 &
      (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_1_mx0w0)) | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_1_mx0w0
      | lfst_exit_PADDING_LOOP_lpi_1_dfm_0_mx0w0));
  assign nl_LOAD_LOOP_i_sva_1_mx0w0 = LOAD_LOOP_i_lpi_1_mx0 + 16'b0000000000000001;
  assign LOAD_LOOP_i_sva_1_mx0w0 = nl_LOAD_LOOP_i_sva_1_mx0w0[15:0];
  assign LOAD_LOOP_LOAD_LOOP_if_and_tmp = (LOAD_LOOP_i_lpi_1_mx0 == (operator_32_false_acc_psp_sva_1[15:0]))
      & (operator_32_false_acc_psp_sva_1[32:16]==17'b00000000000000000);
  assign PADDING_LOOP_equal_tmp_mx1w0 = lfst_exit_PADDING_LOOP_lpi_1_dfm_1_mx0w0
      & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_0_mx0w0);
  assign PADDING_LOOP_equal_tmp_1_mx0w0 = lfst_exit_PADDING_LOOP_lpi_1_dfm_1_mx0w0
      & lfst_exit_PADDING_LOOP_lpi_1_dfm_0_mx0w0;
  assign PADDING_LOOP_for_for_land_2_lpi_1_dfm_mx0w0 = PADDING_LOOP_for_for_aelse_2_acc_itm_9_1
      & PADDING_LOOP_for_for_aelse_1_acc_itm_9_1 & (~(PADDING_LOOP_for_for_aelse_acc_itm_8
      | PADDING_LOOP_for_for_if_acc_itm_8));
  assign nl_operator_16_false_acc_nl = conv_u2u_6_7(LOAD_LOOP_i_sva_1_mx0w0[15:10])
      + 7'b1001111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[6:0];
  assign exit_LOAD_LOOP_lpi_1_dfm_mx1w0 = (~ (readslicef_7_1_6(operator_16_false_acc_nl)))
      | LOAD_LOOP_LOAD_LOOP_if_and_tmp;
  assign PADDING_LOOP_mux_10_nl = MUX_s_1_2_2(lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1,
      lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1_mx0w0, and_5_tmp);
  assign lfst_exit_PADDING_LOOP_lpi_1_dfm_1_mx0w0 = PADDING_LOOP_mux_10_nl & (~ exitL_exit_PADDING_LOOP_lpi_1_dfm_1);
  assign PADDING_LOOP_mux_13_nl = MUX_s_1_2_2(lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0,
      lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0_mx0w0, and_5_tmp);
  assign lfst_exit_PADDING_LOOP_lpi_1_dfm_0_mx0w0 = PADDING_LOOP_mux_13_nl & (~ exitL_exit_PADDING_LOOP_lpi_1_dfm_1);
  assign LOAD_BATCH_LOOP_mux_8_nl = MUX_s_1_2_2(exit_LOAD_BATCH_LOOP_sva_2_mx0w0,
      exit_LOAD_BATCH_LOOP_sva_2, or_tmp_86);
  assign exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_mx0w0 = ((LOAD_BATCH_LOOP_b_4_0_sva_2[4])
      | LOAD_BATCH_LOOP_mux_8_nl) & exit_PADDING_LOOP_lpi_1_dfm_2_mx1 & PADDING_LOOP_equal_tmp_1_mx0w0;
  assign PADDING_LOOP_for_for_and_3_psp_mx1w0 = (~ exit_PADDING_LOOP_for_sva_5) &
      exit_PADDING_LOOP_for_for_lpi_1_dfm_1;
  assign PADDING_LOOP_for_for_and_3_psp_mx1 = MUX_s_1_2_2(PADDING_LOOP_for_for_and_3_psp_mx1w0,
      PADDING_LOOP_for_for_and_3_psp, or_dcpl_39);
  assign PADDING_LOOP_for_and_psp_mx1w0 = (~ exit_PADDING_LOOP_sva_2) & exit_PADDING_LOOP_for_lpi_1_dfm_4;
  assign exit_PADDING_LOOP_for_for_lpi_1_dfm_1 = ~(operator_8_false_3_acc_itm_4_1
      & ((~(PADDING_LOOP_for_for_if_1_equal_tmp & (operator_8_false_1_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_1_acc_tmp[8])));
  assign LOAD_LOOP_mul_1_nl = conv_u2u_24_24(mul_4_cse_lpi_1_dfm * conf_info_crt_lpi_1_dfm_135_128);
  assign LOAD_LOOP_mul_nl = conv_u2u_32_32(LOAD_LOOP_mul_1_nl * conf_info_crt_lpi_1_dfm_71_64);
  assign nl_operator_32_false_acc_psp_sva_1 = conv_u2s_32_33(LOAD_LOOP_mul_nl) +
      33'b111111111111111111111111111111111;
  assign operator_32_false_acc_psp_sva_1 = nl_operator_32_false_acc_psp_sva_1[32:0];
  assign LOAD_BATCH_LOOP_not_17_nl = ~ exitL_exit_LOAD_BATCH_LOOP_sva;
  assign LOAD_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1 = MUX_v_4_2_2(4'b0000, LOAD_BATCH_LOOP_b_4_0_lpi_1_3_0,
      LOAD_BATCH_LOOP_not_17_nl);
  assign nl_LOAD_BATCH_LOOP_b_4_0_sva_2 = conv_u2u_4_5(LOAD_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1)
      + 5'b00001;
  assign LOAD_BATCH_LOOP_b_4_0_sva_2 = nl_LOAD_BATCH_LOOP_b_4_0_sva_2[4:0];
  assign nl_PADDING_LOOP_for_for_aelse_2_acc_1_nl = conv_u2u_8_9({(~ n_w_in_acc_psp_lpi_1_dfm)
      , (~ conf_info_crt_lpi_1_dfm_192)}) + conv_u2u_8_9(pad_lpi_1_dfm) + 9'b000000001;
  assign PADDING_LOOP_for_for_aelse_2_acc_1_nl = nl_PADDING_LOOP_for_for_aelse_2_acc_1_nl[8:0];
  assign nl_PADDING_LOOP_for_for_aelse_2_acc_nl = conv_u2u_9_10(PADDING_LOOP_for_for_aelse_2_acc_1_nl)
      + conv_s2u_9_10({4'b1000 , PADDING_LOOP_for_row_4_0_lpi_1});
  assign PADDING_LOOP_for_for_aelse_2_acc_nl = nl_PADDING_LOOP_for_for_aelse_2_acc_nl[9:0];
  assign PADDING_LOOP_for_for_aelse_2_acc_itm_9_1 = readslicef_10_1_9(PADDING_LOOP_for_for_aelse_2_acc_nl);
  assign nl_PADDING_LOOP_for_for_aelse_1_acc_1_nl = conv_u2u_8_9({(~ n_h_in_acc_psp_lpi_1_dfm)
      , (~ conf_info_crt_lpi_1_dfm_160)}) + conv_u2u_8_9(pad_lpi_1_dfm) + 9'b000000001;
  assign PADDING_LOOP_for_for_aelse_1_acc_1_nl = nl_PADDING_LOOP_for_for_aelse_1_acc_1_nl[8:0];
  assign nl_PADDING_LOOP_for_for_aelse_1_acc_nl = conv_u2u_9_10(PADDING_LOOP_for_for_aelse_1_acc_1_nl)
      + conv_s2u_9_10({4'b1000 , PADDING_LOOP_for_for_col_4_0_lpi_1_dfm_3});
  assign PADDING_LOOP_for_for_aelse_1_acc_nl = nl_PADDING_LOOP_for_for_aelse_1_acc_nl[9:0];
  assign PADDING_LOOP_for_for_aelse_1_acc_itm_9_1 = readslicef_10_1_9(PADDING_LOOP_for_for_aelse_1_acc_nl);
  assign PADDING_LOOP_for_for_col_4_0_lpi_1_dfm_3 = MUX_v_5_2_2(5'b00000, PADDING_LOOP_for_for_col_4_0_lpi_1,
      lfst_exit_PADDING_LOOP_for_1_lpi_1);
  assign nl_PADDING_LOOP_for_for_aelse_acc_nl = ({4'b1000 , PADDING_LOOP_for_for_col_4_0_lpi_1_dfm_3})
      + conv_u2u_8_9(~ pad_lpi_1_dfm) + 9'b000000001;
  assign PADDING_LOOP_for_for_aelse_acc_nl = nl_PADDING_LOOP_for_for_aelse_acc_nl[8:0];
  assign PADDING_LOOP_for_for_aelse_acc_itm_8 = readslicef_9_1_8(PADDING_LOOP_for_for_aelse_acc_nl);
  assign nl_operator_8_false_4_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_231_224)
      + 9'b111111111;
  assign operator_8_false_4_acc_tmp = nl_operator_8_false_4_acc_tmp[8:0];
  assign nl_PADDING_LOOP_acc_tmp = conv_u2u_5_6(PADDING_LOOP_chan_5_0_lpi_1_4_0)
      + 6'b000001;
  assign PADDING_LOOP_acc_tmp = nl_PADDING_LOOP_acc_tmp[5:0];
  assign PADDING_LOOP_if_equal_tmp = PADDING_LOOP_chan_5_0_lpi_1_4_0 == (operator_8_false_3_acc_tmp[4:0]);
  assign exit_PADDING_LOOP_sva_2 = ~((~(PADDING_LOOP_if_equal_tmp & (operator_8_false_3_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_3_acc_tmp[8]));
  assign nl_operator_8_false_3_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_135_128)
      + 9'b111111111;
  assign operator_8_false_3_acc_tmp = nl_operator_8_false_3_acc_tmp[8:0];
  assign nl_operator_8_false_2_acc_nl = conv_u2s_4_5(PADDING_LOOP_for_row_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_2_acc_nl = nl_operator_8_false_2_acc_nl[4:0];
  assign operator_8_false_2_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_2_acc_nl);
  assign nl_PADDING_LOOP_for_row_4_0_sva_2 = PADDING_LOOP_for_row_4_0_lpi_1 + 5'b00001;
  assign PADDING_LOOP_for_row_4_0_sva_2 = nl_PADDING_LOOP_for_row_4_0_sva_2[4:0];
  assign PADDING_LOOP_for_if_equal_tmp = PADDING_LOOP_for_row_4_0_lpi_1 == (operator_8_false_2_acc_tmp[4:0]);
  assign exit_PADDING_LOOP_for_sva_5 = ~((~(PADDING_LOOP_for_if_equal_tmp & (operator_8_false_2_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_2_acc_tmp[8]));
  assign nl_operator_8_false_2_acc_tmp = conv_u2s_8_9({n_w_in_acc_psp_lpi_1_dfm ,
      conf_info_crt_lpi_1_dfm_192}) + 9'b111111111;
  assign operator_8_false_2_acc_tmp = nl_operator_8_false_2_acc_tmp[8:0];
  assign nl_operator_8_false_3_acc_nl = conv_u2s_4_5(PADDING_LOOP_for_for_col_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_3_acc_nl = nl_operator_8_false_3_acc_nl[4:0];
  assign operator_8_false_3_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_3_acc_nl);
  assign nl_PADDING_LOOP_for_for_col_4_0_sva_2 = PADDING_LOOP_for_for_col_4_0_lpi_1_dfm_3
      + 5'b00001;
  assign PADDING_LOOP_for_for_col_4_0_sva_2 = nl_PADDING_LOOP_for_for_col_4_0_sva_2[4:0];
  assign PADDING_LOOP_for_mux_1_nl = MUX_s_1_2_2(exit_PADDING_LOOP_for_lpi_1_dfm_1_mx0w0,
      exit_PADDING_LOOP_for_lpi_1_dfm_1, and_197_cse);
  assign exit_PADDING_LOOP_for_lpi_1_dfm_4 = PADDING_LOOP_for_mux_1_nl & exit_PADDING_LOOP_for_for_lpi_1_dfm_1;
  assign PADDING_LOOP_for_for_if_1_equal_tmp = PADDING_LOOP_for_for_col_4_0_lpi_1_dfm_3
      == (operator_8_false_1_acc_tmp[4:0]);
  assign nl_operator_8_false_1_acc_tmp = conv_u2s_8_9({n_h_in_acc_psp_lpi_1_dfm ,
      conf_info_crt_lpi_1_dfm_160}) + 9'b111111111;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[8:0];
  assign nl_PADDING_LOOP_for_for_if_acc_nl = ({4'b1000 , PADDING_LOOP_for_row_4_0_lpi_1})
      + conv_u2u_8_9(~ pad_lpi_1_dfm) + 9'b000000001;
  assign PADDING_LOOP_for_for_if_acc_nl = nl_PADDING_LOOP_for_for_if_acc_nl[8:0];
  assign PADDING_LOOP_for_for_if_acc_itm_8 = readslicef_9_1_8(PADDING_LOOP_for_for_if_acc_nl);
  assign PADDING_LOOP_and_2_ssc_1 = dma_read_ctrl_rsci_irdy_mxwt & PADDING_LOOP_or_tmp_1;
  assign nl_ac_int_cctor_8_sva_1 = z_out_1 + z_out_2;
  assign ac_int_cctor_8_sva_1 = nl_ac_int_cctor_8_sva_1[15:0];
  assign mul_4_cse_sva_1 = conv_u2u_16_16((conf_info_rsci_idat_mxwt[31:24]) * (conf_info_rsci_idat_mxwt[31:24]));
  assign operator_43_true_and_nl = (pad_acc_psp_sva_1[16]) & (pad_acc_psp_sva_1[0]);
  assign nl_operator_43_true_operator_43_true_acc_nl = (pad_acc_psp_sva_1[8:1]) +
      conv_u2s_1_8(operator_43_true_and_nl);
  assign operator_43_true_operator_43_true_acc_nl = nl_operator_43_true_operator_43_true_acc_nl[7:0];
  assign nl_pad_sva_1 = $signed(operator_43_true_operator_43_true_acc_nl) * $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[15:8]));
  assign pad_sva_1 = nl_pad_sva_1[7:0];
  assign exitL_exit_PADDING_LOOP_lpi_1_dfm_1 = exitL_exit_PADDING_LOOP_lpi_1_mx0
      | exit_LOAD_BATCH_LOOP_lpi_1_dfm_3 | exitL_exit_LOAD_BATCH_LOOP_sva;
  assign and_7_tmp = (conf_info_rsci_bawt | (~ LOAD_BATCH_LOOP_asn_itm)) & (dma_read_ctrl_rsci_bawt
      | (~(((lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0 & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1))
      | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 | lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0)))
      & main_stage_v_1))) & (dma_read_chnl_rsci_bawt | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1
      & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0) & main_stage_v_1))) & or_10_cse_1
      & or_11_cse_1 & or_12_cse_1 & or_13_cse_1 & or_4_cse_1 & or_5_cse_1 & or_6_cse_1
      & or_cse_1;
  assign or_10_cse_1 = dma_read_chnl_rsci_bawt | (~(PADDING_LOOP_for_for_land_2_lpi_1_dfm_st_1
      & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0
      & main_stage_v_1));
  assign or_11_cse_1 = plm_filters_rsc_req_obj_bawt | nand_21_cse_1;
  assign or_12_cse_1 = plm_inputs_rsc_req_obj_bawt | nand_21_cse_1;
  assign or_13_cse_1 = plm_filters_rsci_bawt | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1
      & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0) & main_stage_v_2));
  assign or_4_cse_1 = plm_inputs_rsci_bawt | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1
      & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0 & main_stage_v_2));
  assign or_5_cse_1 = plm_filters_rsc_rls_obj_bawt | nand_9_cse_1;
  assign or_6_cse_1 = plm_inputs_rsc_rls_obj_bawt | nand_9_cse_1;
  assign or_cse_1 = done_rsci_bawt | (~(exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_3 & main_stage_v_3));
  assign nand_21_cse_1 = ~(exit_LOAD_CTRL_LOOP_sva_st_1 & PADDING_LOOP_or_cse_1 &
      main_stage_v_2);
  assign PADDING_LOOP_or_cse_1 = (lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0 & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1))
      | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1 | lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0));
  assign nand_5_cse_1 = ~(exit_LOAD_CTRL_LOOP_sva_st_1 & PADDING_LOOP_or_cse_1);
  assign nand_9_cse_1 = ~(exit_PADDING_LOOP_lpi_1_dfm_2_st_2 & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1
      & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0 & main_stage_v_2);
  assign PADDING_LOOP_and_8_m1c_1 = (~ exit_PADDING_LOOP_for_lpi_1_dfm_4) & PADDING_LOOP_equal_tmp_1_mx0w0;
  assign nl_pad_acc_2_nl = ({1'b1 , (~ (conf_info_rsci_idat_mxwt[55:48]))}) + conv_u2s_8_9(conf_info_rsci_idat_mxwt[31:24])
      + 9'b000000001;
  assign pad_acc_2_nl = nl_pad_acc_2_nl[8:0];
  assign nl_operator_8_false_acc_nl = conv_u2s_8_9(conf_info_rsci_idat_mxwt[55:48])
      + 9'b111111111;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[8:0];
  assign nl_pad_mul_nl = $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[7:0])) * $signed(operator_8_false_acc_nl);
  assign pad_mul_nl = nl_pad_mul_nl[16:0];
  assign nl_pad_acc_psp_sva_1 = conv_s2s_9_17(pad_acc_2_nl) + pad_mul_nl;
  assign pad_acc_psp_sva_1 = nl_pad_acc_psp_sva_1[16:0];
  assign and_5_tmp = main_stage_v_1 & (dma_read_ctrl_rsci_bawt | lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1)
      & (dma_read_chnl_rsci_bawt | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 & (~
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0)))) & or_10_cse_1 & or_11_cse_1 & or_12_cse_1
      & or_13_cse_1 & or_4_cse_1 & or_5_cse_1 & or_6_cse_1 & or_cse_1;
  assign and_3_tmp = main_stage_v_2 & (plm_filters_rsc_req_obj_bawt | nand_5_cse_1)
      & (plm_inputs_rsc_req_obj_bawt | nand_5_cse_1) & (plm_filters_rsci_bawt | (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1
      & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0)))) & or_4_cse_1 & or_5_cse_1
      & or_6_cse_1 & or_cse_1;
  assign or_tmp_3 = lfst_exit_PADDING_LOOP_lpi_1_dfm_2_1_0 | PADDING_LOOP_equal_tmp_1_1;
  assign or_tmp_10 = exitL_exit_LOAD_BATCH_LOOP_sva | exit_LOAD_BATCH_LOOP_lpi_1_dfm_3;
  assign or_tmp_18 = (~((~ PADDING_LOOP_if_equal_tmp) | (operator_8_false_3_acc_tmp[8:5]!=4'b0000)))
      | (PADDING_LOOP_acc_tmp[5]);
  assign or_62_cse = (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1) | (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0)
      | exitL_exit_PADDING_LOOP_lpi_1;
  assign or_73_cse = (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1) | exitL_exit_PADDING_LOOP_lpi_1;
  assign or_tmp_64 = or_tmp_10 | mux_70_cse;
  assign or_115_nl = or_62_cse | (~ or_tmp_18);
  assign nand_66_nl = ~(lfst_exit_PADDING_LOOP_lpi_1_dfm_2_1_0 & or_tmp_18);
  assign nand_67_nl = ~(lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0 & or_tmp_18);
  assign mux_18_nl = MUX_s_1_2_2(nand_66_nl, nand_67_nl, PADDING_LOOP_equal_tmp_1_1);
  assign or_50_nl = PADDING_LOOP_or_tmp_1 | mux_18_nl;
  assign mux_tmp_65 = MUX_s_1_2_2(or_115_nl, or_50_nl, and_5_tmp);
  assign or_118_nl = or_tmp_10 | mux_tmp_65;
  assign or_116_nl = (~ PADDING_LOOP_for_for_if_1_equal_tmp) | (operator_8_false_1_acc_tmp[8:5]!=4'b0000)
      | exitL_exit_LOAD_BATCH_LOOP_sva | exit_LOAD_BATCH_LOOP_lpi_1_dfm_3 | mux_tmp_65;
  assign mux_66_nl = MUX_s_1_2_2(or_118_nl, or_116_nl, operator_8_false_3_acc_itm_4_1);
  assign or_tmp_86 = and_193_cse | mux_66_nl;
  assign and_dcpl_1 = and_7_tmp & LOAD_BATCH_LOOP_asn_itm;
  assign or_126_nl = (~ PADDING_LOOP_for_for_if_1_equal_tmp) | (operator_8_false_1_acc_tmp[8:5]!=4'b0000)
      | mux_tmp_65;
  assign mux_68_nl = MUX_s_1_2_2(mux_tmp_65, or_126_nl, operator_8_false_3_acc_itm_4_1);
  assign or_tmp_92 = and_193_cse | mux_68_nl;
  assign nor_40_nl = ~(PADDING_LOOP_or_tmp_1 | (~ PADDING_LOOP_equal_tmp_1_1) | lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0);
  assign not_tmp_61 = MUX_s_1_2_2(exitL_exit_PADDING_LOOP_lpi_1, nor_40_nl, and_5_tmp);
  assign and_dcpl_4 = (~ exitL_exit_LOAD_BATCH_LOOP_sva) & and_7_tmp;
  assign and_dcpl_6 = ~(exit_LOAD_BATCH_LOOP_lpi_1_dfm_3 | exitL_exit_LOAD_BATCH_LOOP_sva);
  assign and_dcpl_7 = and_dcpl_6 & and_7_tmp;
  assign or_tmp_109 = lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 | (~ dma_read_ctrl_rsci_irdy_mxwt);
  assign mux_75_nl = MUX_s_1_2_2(or_42_cse, (~ or_tmp_109), PADDING_LOOP_or_tmp_1);
  assign mux_tmp_76 = MUX_s_1_2_2((~ or_73_cse), mux_75_nl, and_5_tmp);
  assign and_dcpl_15 = and_3_tmp & (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1) &
      exit_LOAD_CTRL_LOOP_sva_st_1;
  assign and_dcpl_16 = and_dcpl_15 & (or_tmp_109 | (~ and_5_tmp));
  assign and_dcpl_19 = lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0 & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1;
  assign and_dcpl_22 = and_3_tmp & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1;
  assign and_dcpl_26 = main_stage_v_3 & done_rsci_bawt & exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_3;
  assign and_dcpl_27 = and_dcpl_26 & (~(and_3_tmp & exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_2));
  assign or_162_cse = (~ PADDING_LOOP_for_for_aelse_2_acc_itm_9_1) | (~ PADDING_LOOP_for_for_aelse_1_acc_itm_9_1)
      | PADDING_LOOP_for_for_aelse_acc_itm_8 | PADDING_LOOP_for_for_if_acc_itm_8;
  assign mux_13_nl = MUX_s_1_2_2(or_42_cse, dma_read_ctrl_rsci_irdy_mxwt, PADDING_LOOP_or_tmp_1);
  assign mux_81_nl = MUX_s_1_2_2((~ or_73_cse), mux_13_nl, and_5_tmp);
  assign mux_78_nl = MUX_s_1_2_2((~ or_tmp_3), dma_read_ctrl_rsci_irdy_mxwt, PADDING_LOOP_or_tmp_1);
  assign mux_79_nl = MUX_s_1_2_2((~ or_38_cse), mux_78_nl, and_5_tmp);
  assign mux_82_nl = MUX_s_1_2_2(mux_81_nl, mux_79_nl, or_162_cse);
  assign and_dcpl_29 = mux_82_nl & and_dcpl_7;
  assign and_dcpl_30 = lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 & and_5_tmp;
  assign or_dcpl_18 = (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0) | PADDING_LOOP_for_for_land_2_lpi_1_dfm_st_1;
  assign or_dcpl_19 = or_tmp_10 | (~ and_7_tmp);
  assign mux_tmp_85 = MUX_s_1_2_2(dma_read_ctrl_rsci_irdy_mxwt, or_dcpl_18, lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1);
  assign not_tmp_85 = ~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 & or_dcpl_18);
  assign or_dcpl_23 = lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0 | (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1)
      | (~ and_5_tmp);
  assign or_dcpl_25 = ~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0 & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1
      & and_5_tmp);
  assign or_196_nl = (~ PADDING_LOOP_for_for_if_1_equal_tmp) | (operator_8_false_1_acc_tmp[8:5]!=4'b0000)
      | mux_70_cse;
  assign mux_tmp_95 = MUX_s_1_2_2(mux_70_cse, or_196_nl, operator_8_false_3_acc_itm_4_1);
  assign and_dcpl_54 = (~ mux_70_cse) & and_dcpl_7;
  assign or_205_nl = PADDING_LOOP_or_tmp_1 | (~ or_tmp_3);
  assign mux_96_nl = MUX_s_1_2_2((~ lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0), or_205_nl,
      and_5_tmp);
  assign or_dcpl_39 = mux_96_nl | or_tmp_10;
  assign nor_24_cse = ~((~((~ LOAD_BATCH_LOOP_if_1_equal_tmp) | (operator_8_false_4_acc_tmp[8:4]!=5'b00000)))
      | (LOAD_BATCH_LOOP_b_4_0_sva_2[4]));
  assign or_tmp_137 = (nor_24_cse | or_tmp_92 | or_tmp_10 | (~ and_7_tmp)) & and_dcpl_1
      & (fsm_output[1]);
  assign or_tmp_152 = (~ lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1) & and_5_tmp & (fsm_output[1]);
  assign and_165_cse = or_tmp_64 & and_7_tmp & (fsm_output[1]);
  assign nor_18_nl = ~(lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1 | exitL_exit_PADDING_LOOP_lpi_1);
  assign and_194_nl = PADDING_LOOP_or_tmp_1 & or_tmp_109;
  assign mux_74_nl = MUX_s_1_2_2(nor_18_nl, and_194_nl, and_5_tmp);
  assign dma_read_ctrl_rsci_idat_15_0_mx0c1 = mux_74_nl & and_dcpl_7;
  assign dma_read_ctrl_rsci_idat_47_32_mx0c1 = ((~ mux_tmp_76) | exit_LOAD_BATCH_LOOP_lpi_1_dfm_3)
      & and_dcpl_4;
  assign main_stage_v_3_mx0c1 = (done_rsci_bawt | (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_3))
      & main_stage_v_3 & (~ and_3_tmp);
  assign main_stage_v_2_mx0c1 = and_3_tmp & (~ and_5_tmp) & (fsm_output[1]);
  assign main_stage_v_1_mx0c1 = and_5_tmp & (~ and_7_tmp) & (fsm_output[1]);
  assign exit_PADDING_LOOP_lpi_1_dfm_2_st_1_mx0c1 = and_165_cse | ((mux_70_cse |
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_3) & and_dcpl_4);
  assign plm_inputs_rsci_d_d = PADDING_LOOP_for_for_mux_rmff;
  assign plm_inputs_rsci_wadr_d = PADDING_LOOP_for_for_index_in_mux_rmff;
  assign plm_inputs_rsci_we_d_pff = plm_inputs_rsci_we_d_iff;
  assign plm_filters_rsci_d_d = LOAD_LOOP_data_ac_mux_rmff;
  assign plm_filters_rsci_wadr_d = LOAD_LOOP_i_mux_rmff;
  assign plm_filters_rsci_we_d_pff = plm_filters_rsci_we_d_iff;
  assign and_dcpl_58 = PADDING_LOOP_equal_tmp_1_mx0w0 & exit_PADDING_LOOP_for_lpi_1_dfm_4;
  assign and_223_cse = exitL_exit_LOAD_BATCH_LOOP_sva & (fsm_output[1]);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (((~(nor_24_cse | or_tmp_86)) & and_7_tmp) | (fsm_output[0])
        | or_tmp_137) ) begin
      reg_conf_info_rsci_iswt0_cse <= ~ or_tmp_137;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exitL_exit_LOAD_BATCH_LOOP_sva <= 1'b1;
      PADDING_LOOP_or_tmp_1 <= 1'b0;
      PADDING_LOOP_equal_tmp_1_1 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0 <= 1'b0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( LOAD_BATCH_LOOP_and_cse ) begin
      exitL_exit_LOAD_BATCH_LOOP_sva <= exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_mx0w0;
      PADDING_LOOP_or_tmp_1 <= PADDING_LOOP_or_tmp_mx0w0;
      PADDING_LOOP_equal_tmp_1_1 <= PADDING_LOOP_equal_tmp_1_mx0w0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_3_1_0 <= ~ exit_PADDING_LOOP_lpi_1_dfm_2_mx1;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 <= lfst_exit_PADDING_LOOP_lpi_1_dfm_1_mx0w0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0 <= lfst_exit_PADDING_LOOP_lpi_1_dfm_0_mx0w0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_3 <= exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_idat_15_0 <= 16'b0000000000000000;
    end
    else if ( core_wen & (((not_tmp_61 | or_tmp_10) & and_7_tmp & (fsm_output[1]))
        | ((not_tmp_61 | exit_LOAD_BATCH_LOOP_lpi_1_dfm_3) & and_dcpl_4) | dma_read_ctrl_rsci_idat_15_0_mx0c1)
        ) begin
      dma_read_ctrl_rsci_idat_15_0 <= MUX_v_16_2_2(LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm_mx0w0,
          LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm, dma_read_ctrl_rsci_idat_15_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( core_wen & ((exitL_exit_LOAD_BATCH_LOOP_sva & and_7_tmp & (fsm_output[1]))
        | dma_read_ctrl_rsci_idat_47_32_mx0c1) ) begin
      dma_read_ctrl_rsci_idat_47_32 <= MUX_v_16_2_2(ac_int_cctor_8_sva_1, ac_int_cctor_8_lpi_1_dfm,
          dma_read_ctrl_rsci_idat_47_32_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_filters_rsc_req_obj_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (((~ or_tmp_109) & and_5_tmp & (fsm_output[1])) | and_dcpl_16)
        ) begin
      reg_plm_filters_rsc_req_obj_iswt0_cse <= ~ and_dcpl_16;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_filters_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_dma_read_ctrl_rsci_ivld_core_psct_cse <= 1'b0;
      reg_plm_filters_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= 1'b0;
      reg_plm_inputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= 1'b0;
      plm_filters_rsci_wadr_d_reg <= 16'b0000000000000000;
      plm_filters_rsci_d_d_reg <= 32'b00000000000000000000000000000000;
      plm_inputs_rsci_wadr_d_reg <= 14'b00000000000000;
      plm_inputs_rsci_d_d_reg <= 32'b00000000000000000000000000000000;
      LOAD_LOOP_i_lpi_1 <= 16'b0000000000000000;
      ac_int_cctor_8_lpi_1_dfm <= 16'b0000000000000000;
      exitL_exit_PADDING_LOOP_lpi_1 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_plm_filters_rsc_rls_obj_ld_core_psct_cse <= and_dcpl_19 & and_5_tmp & exit_PADDING_LOOP_lpi_1_dfm_2_st_1;
      reg_dma_read_ctrl_rsci_ivld_core_psct_cse <= ((~ mux_tmp_76) | or_tmp_10) &
          and_7_tmp & (fsm_output[1]);
      reg_plm_filters_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= and_58_rmff;
      reg_plm_inputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= and_60_rmff;
      plm_filters_rsci_wadr_d_reg <= LOAD_LOOP_i_mux_rmff;
      plm_filters_rsci_d_d_reg <= LOAD_LOOP_data_ac_mux_rmff;
      plm_inputs_rsci_wadr_d_reg <= PADDING_LOOP_for_for_index_in_mux_rmff;
      plm_inputs_rsci_d_d_reg <= PADDING_LOOP_for_for_mux_rmff;
      LOAD_LOOP_i_lpi_1 <= LOAD_LOOP_i_lpi_1_mx0;
      ac_int_cctor_8_lpi_1_dfm <= ac_int_cctor_8_lpi_1_dfm_mx0;
      exitL_exit_PADDING_LOOP_lpi_1 <= exitL_exit_PADDING_LOOP_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_done_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((and_3_tmp & exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_2) | and_dcpl_27)
        ) begin
      reg_done_rsci_ivld_core_psct_cse <= ~ and_dcpl_27;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_read_chnl_rsci_irdy_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (mux_91_nl | and_dcpl_29) ) begin
      reg_dma_read_chnl_rsci_irdy_core_psct_cse <= (~((mux_83_nl | or_dcpl_19) &
          or_dcpl_18 & and_dcpl_30)) | and_dcpl_29;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_asn_itm <= 1'b1;
    end
    else if ( core_wen & and_115_cse ) begin
      LOAD_BATCH_LOOP_asn_itm <= exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & ((and_3_tmp & (fsm_output[1])) | main_stage_v_3_mx0c1) )
        begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_3 <= 1'b0;
    end
    else if ( core_wen & (~((~ and_3_tmp) | (fsm_output[0]))) ) begin
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_3 <= exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & ((and_5_tmp & (fsm_output[1])) | main_stage_v_2_mx0c1) )
        begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_CTRL_LOOP_sva_st_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_152 | and_dcpl_30) ) begin
      exit_LOAD_CTRL_LOOP_sva_st_1 <= MUX_s_1_2_2(dma_read_ctrl_rsci_irdy_mxwt, exit_LOAD_CTRL_LOOP_sva_st,
          and_dcpl_30);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_PADDING_LOOP_lpi_1_dfm_2_st_2 <= 1'b0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_2 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0 <= 1'b0;
    end
    else if ( PADDING_LOOP_and_cse ) begin
      exit_PADDING_LOOP_lpi_1_dfm_2_st_2 <= exit_PADDING_LOOP_lpi_1_dfm_2_st_1;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_3_st_2 <= exit_LOAD_BATCH_LOOP_lpi_1_dfm_3;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_1 <= lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_st_2_0 <= lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1 <= lfst_exit_PADDING_LOOP_lpi_1_dfm_4_1_mx0w0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0 <= lfst_exit_PADDING_LOOP_lpi_1_dfm_4_0_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm <= 16'b0000000000000000;
    end
    else if ( core_wen & (~(mux_92_nl & and_dcpl_6)) & and_7_tmp ) begin
      LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm <= LOAD_BATCH_LOOP_dma_read_info_index_15_0_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      mul_4_cse_lpi_1_dfm <= 16'b0000000000000000;
      conf_info_crt_lpi_1_dfm_135_128 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_71_64 <= 8'b00000000;
      n_w_in_acc_psp_lpi_1_dfm <= 7'b0000000;
      conf_info_crt_lpi_1_dfm_192 <= 1'b0;
      pad_lpi_1_dfm <= 8'b00000000;
      n_h_in_acc_psp_lpi_1_dfm <= 7'b0000000;
      conf_info_crt_lpi_1_dfm_160 <= 1'b0;
      conf_info_crt_lpi_1_dfm_231_224 <= 8'b00000000;
    end
    else if ( and_234_cse ) begin
      mul_4_cse_lpi_1_dfm <= mul_4_cse_sva_1;
      conf_info_crt_lpi_1_dfm_135_128 <= conf_info_rsci_idat_mxwt[39:32];
      conf_info_crt_lpi_1_dfm_71_64 <= conf_info_rsci_idat_mxwt[23:16];
      n_w_in_acc_psp_lpi_1_dfm <= nl_n_w_in_acc_psp_lpi_1_dfm[6:0];
      conf_info_crt_lpi_1_dfm_192 <= conf_info_rsci_idat_mxwt[48];
      pad_lpi_1_dfm <= pad_sva_1;
      n_h_in_acc_psp_lpi_1_dfm <= nl_n_h_in_acc_psp_lpi_1_dfm[6:0];
      conf_info_crt_lpi_1_dfm_160 <= conf_info_rsci_idat_mxwt[40];
      conf_info_crt_lpi_1_dfm_231_224 <= conf_info_rsci_idat_mxwt[63:56];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_BATCH_LOOP_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~(or_tmp_92 | or_dcpl_19)) ) begin
      exit_LOAD_BATCH_LOOP_sva_2 <= exit_LOAD_BATCH_LOOP_sva_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_exit_PADDING_LOOP_lpi_1_dfm_2_cse <= 1'b0;
      PADDING_LOOP_for_for_and_3_psp <= 1'b0;
      PADDING_LOOP_for_and_psp <= 1'b0;
      PADDING_LOOP_for_for_land_2_lpi_1_dfm_st <= 1'b0;
    end
    else if ( PADDING_LOOP_and_31_cse ) begin
      reg_exit_PADDING_LOOP_lpi_1_dfm_2_cse <= exit_PADDING_LOOP_lpi_1_dfm_2_mx1w0;
      PADDING_LOOP_for_for_and_3_psp <= PADDING_LOOP_for_for_and_3_psp_mx1w0;
      PADDING_LOOP_for_and_psp <= PADDING_LOOP_for_and_psp_mx1w0;
      PADDING_LOOP_for_for_land_2_lpi_1_dfm_st <= PADDING_LOOP_for_for_land_2_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_for_row_4_0_lpi_1 <= 5'b00000;
    end
    else if ( core_wen & (~((and_dcpl_58 & exit_PADDING_LOOP_lpi_1_dfm_mx0w0 & (~
        PADDING_LOOP_for_for_and_3_psp_mx1w0)) | ((~ PADDING_LOOP_for_for_and_3_psp_mx1)
        & PADDING_LOOP_and_8_m1c_1) | (~ and_7_tmp) | PADDING_LOOP_or_tmp_mx0w0))
        ) begin
      PADDING_LOOP_for_row_4_0_lpi_1 <= MUX_v_5_2_2((signext_5_1(PADDING_LOOP_for_row_PADDING_LOOP_for_row_PADDING_LOOP_for_row_mux_nl)),
          PADDING_LOOP_for_row_4_0_sva_2, and_217_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_PADDING_LOOP_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(and_193_cse | mux_tmp_95 | or_dcpl_19)) ) begin
      exit_PADDING_LOOP_lpi_1_dfm <= exit_PADDING_LOOP_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_chan_5_0_lpi_1_4_0 <= 5'b00000;
    end
    else if ( core_wen & ((PADDING_LOOP_equal_tmp_mx1w0 & and_7_tmp) | PADDING_LOOP_and_7_rgt)
        ) begin
      PADDING_LOOP_chan_5_0_lpi_1_4_0 <= MUX_v_5_2_2((signext_5_1(~ exit_LOAD_LOOP_lpi_1_dfm_mx1w0)),
          (PADDING_LOOP_acc_tmp[4:0]), PADDING_LOOP_and_7_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_PADDING_LOOP_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(mux_tmp_95 | or_dcpl_19)) ) begin
      exit_PADDING_LOOP_for_lpi_1_dfm_1 <= exit_PADDING_LOOP_for_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_for_for_col_4_0_lpi_1 <= 5'b00000;
    end
    else if ( core_wen & (((~ exit_PADDING_LOOP_for_for_lpi_1_dfm_1) & PADDING_LOOP_equal_tmp_1_mx0w0
        & and_7_tmp) | PADDING_LOOP_and_11_rgt) ) begin
      PADDING_LOOP_for_for_col_4_0_lpi_1 <= MUX_v_5_2_2(PADDING_LOOP_for_for_col_4_0_sva_2,
          ({{4{exit_PADDING_LOOP_for_lpi_1_dfm_1_mx0w0}}, exit_PADDING_LOOP_for_lpi_1_dfm_1_mx0w0}),
          PADDING_LOOP_and_11_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_PADDING_LOOP_for_1_lpi_1 <= 1'b0;
    end
    else if ( core_wen & (PADDING_LOOP_equal_tmp_mx1w0 | PADDING_LOOP_equal_tmp_1_mx0w0)
        & and_7_tmp ) begin
      lfst_exit_PADDING_LOOP_for_1_lpi_1 <= MUX_s_1_2_2(LOAD_LOOP_LOAD_LOOP_and_2_nl,
          (~ exit_PADDING_LOOP_for_lpi_1_dfm_4), PADDING_LOOP_equal_tmp_1_mx0w0);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_BATCH_LOOP_b_4_0_lpi_1_3_0 <= 4'b0000;
    end
    else if ( core_wen & (((~ or_tmp_92) & and_dcpl_7) | and_73_rgt) ) begin
      LOAD_BATCH_LOOP_b_4_0_lpi_1_3_0 <= MUX_v_4_2_2((LOAD_BATCH_LOOP_b_4_0_sva_2[3:0]),
          LOAD_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1, and_73_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (and_115_cse | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_i_sva_1_1 <= 16'b0000000000000000;
      PADDING_LOOP_for_for_land_2_lpi_1_dfm_1 <= 1'b0;
      PADDING_LOOP_for_for_index_in_acc_itm_1 <= 14'b00000000000000;
    end
    else if ( LOAD_LOOP_i_and_cse ) begin
      LOAD_LOOP_i_sva_1_1 <= LOAD_LOOP_i_sva_1_mx0w0;
      PADDING_LOOP_for_for_land_2_lpi_1_dfm_1 <= PADDING_LOOP_for_for_land_2_lpi_1_dfm_mx0w0;
      PADDING_LOOP_for_for_index_in_acc_itm_1 <= nl_PADDING_LOOP_for_for_index_in_acc_itm_1[13:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_LOOP_sva_1 <= 1'b0;
      PADDING_LOOP_equal_tmp_1 <= 1'b0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_2_1_0 <= 1'b0;
    end
    else if ( LOAD_LOOP_and_cse ) begin
      exit_LOAD_LOOP_sva_1 <= LOAD_LOOP_LOAD_LOOP_if_and_tmp;
      PADDING_LOOP_equal_tmp_1 <= PADDING_LOOP_equal_tmp_mx1w0;
      lfst_exit_PADDING_LOOP_lpi_1_dfm_2_1_0 <= exit_LOAD_LOOP_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_PADDING_LOOP_lpi_1_dfm_2_st_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_54 | exit_PADDING_LOOP_lpi_1_dfm_2_st_1_mx0c1)
        ) begin
      exit_PADDING_LOOP_lpi_1_dfm_2_st_1 <= MUX_s_1_2_2(exit_PADDING_LOOP_lpi_1_dfm_2_mx1w0,
          reg_exit_PADDING_LOOP_lpi_1_dfm_2_cse, exit_PADDING_LOOP_lpi_1_dfm_2_st_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      PADDING_LOOP_for_for_land_2_lpi_1_dfm_st_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_54 | and_165_cse) ) begin
      PADDING_LOOP_for_for_land_2_lpi_1_dfm_st_1 <= MUX_s_1_2_2(PADDING_LOOP_for_for_land_2_lpi_1_dfm_mx0w0,
          PADDING_LOOP_for_for_land_2_lpi_1_dfm_st, and_165_cse);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_CTRL_LOOP_sva_st <= 1'b0;
    end
    else if ( core_wen & (~(lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 | (~ and_5_tmp)))
        ) begin
      exit_LOAD_CTRL_LOOP_sva_st <= dma_read_ctrl_rsci_irdy_mxwt;
    end
  end
  assign mux_83_nl = MUX_s_1_2_2((~ or_42_cse), or_tmp_3, or_162_cse);
  assign and_53_nl = and_5_tmp & lfst_exit_PADDING_LOOP_lpi_1_dfm_st_1_1 & or_dcpl_18;
  assign nand_49_nl = ~(PADDING_LOOP_nor_cse & not_tmp_85);
  assign mux_88_nl = MUX_s_1_2_2(nand_49_nl, mux_tmp_85, PADDING_LOOP_or_tmp_1);
  assign mux_89_nl = MUX_s_1_2_2((~ or_73_cse), mux_88_nl, and_5_tmp);
  assign nand_48_nl = ~(or_tmp_3 & not_tmp_85);
  assign mux_86_nl = MUX_s_1_2_2(nand_48_nl, mux_tmp_85, PADDING_LOOP_or_tmp_1);
  assign mux_87_nl = MUX_s_1_2_2((~ or_38_cse), mux_86_nl, and_5_tmp);
  assign mux_90_nl = MUX_s_1_2_2(mux_89_nl, mux_87_nl, or_162_cse);
  assign nor_13_nl = ~(exitL_exit_LOAD_BATCH_LOOP_sva | exit_LOAD_BATCH_LOOP_lpi_1_dfm_3
      | (~ and_7_tmp));
  assign mux_91_nl = MUX_s_1_2_2(and_53_nl, mux_90_nl, nor_13_nl);
  assign mux_92_nl = MUX_s_1_2_2((~ exitL_exit_PADDING_LOOP_lpi_1), PADDING_LOOP_or_tmp_1,
      and_5_tmp);
  assign nl_n_w_in_acc_psp_lpi_1_dfm  = (conf_info_rsci_idat_mxwt[55:49]) + (pad_sva_1[6:0]);
  assign nl_n_h_in_acc_psp_lpi_1_dfm  = (conf_info_rsci_idat_mxwt[47:41]) + (pad_sva_1[6:0]);
  assign PADDING_LOOP_and_9_nl = exit_PADDING_LOOP_for_lpi_1_dfm_4 & PADDING_LOOP_equal_tmp_1_mx0w0
      & and_7_tmp;
  assign PADDING_LOOP_for_row_PADDING_LOOP_for_row_PADDING_LOOP_for_row_mux_nl =
      MUX_s_1_2_2((~ exit_LOAD_LOOP_lpi_1_dfm_mx1w0), exit_PADDING_LOOP_lpi_1_dfm_mx0w0,
      PADDING_LOOP_and_9_nl);
  assign and_217_nl = ((and_dcpl_58 & exit_PADDING_LOOP_lpi_1_dfm_mx0w0 & PADDING_LOOP_for_for_and_3_psp_mx1w0)
      | (PADDING_LOOP_for_for_and_3_psp_mx1 & PADDING_LOOP_and_8_m1c_1)) & and_7_tmp;
  assign LOAD_LOOP_LOAD_LOOP_and_2_nl = lfst_exit_PADDING_LOOP_for_1_lpi_1 & (~ exit_LOAD_LOOP_lpi_1_dfm_mx1w0);
  assign nl_PADDING_LOOP_for_for_index_in_acc_2_nl = (z_out[12:0]) + conv_u2u_5_13(PADDING_LOOP_for_for_col_4_0_lpi_1_dfm_3);
  assign PADDING_LOOP_for_for_index_in_acc_2_nl = nl_PADDING_LOOP_for_for_index_in_acc_2_nl[12:0];
  assign nl_PADDING_LOOP_for_for_index_in_acc_itm_1  = conv_u2u_13_14(PADDING_LOOP_for_for_index_in_acc_2_nl)
      + (z_out_2[13:0]);
  assign PADDING_LOOP_for_for_index_in_mux_8_nl = MUX_v_8_2_2(({n_h_in_acc_psp_lpi_1_dfm
      , conf_info_crt_lpi_1_dfm_160}), (conf_info_rsci_idat_mxwt[39:32]), and_223_cse);
  assign PADDING_LOOP_for_for_index_in_mux_9_nl = MUX_v_16_2_2(({11'b00000000000
      , PADDING_LOOP_for_row_4_0_lpi_1}), mul_4_cse_sva_1, and_223_cse);
  assign nl_z_out = PADDING_LOOP_for_for_index_in_mux_8_nl * PADDING_LOOP_for_for_index_in_mux_9_nl;
  assign z_out = nl_z_out[15:0];
  assign PADDING_LOOP_for_for_index_in_mux_10_nl = MUX_v_8_2_2(({n_w_in_acc_psp_lpi_1_dfm
      , conf_info_crt_lpi_1_dfm_192}), (conf_info_rsci_idat_mxwt[39:32]), and_223_cse);
  assign mul_6_nl = conv_u2u_16_16((conf_info_rsci_idat_mxwt[55:48]) * (conf_info_rsci_idat_mxwt[47:40]));
  assign PADDING_LOOP_for_for_index_in_mux_11_nl = MUX_v_16_2_2(({11'b00000000000
      , PADDING_LOOP_chan_5_0_lpi_1_4_0}), mul_6_nl, and_223_cse);
  assign nl_z_out_1 = PADDING_LOOP_for_for_index_in_mux_10_nl * PADDING_LOOP_for_for_index_in_mux_11_nl;
  assign z_out_1 = nl_z_out_1[15:0];
  assign PADDING_LOOP_for_for_index_in_mux_12_nl = MUX_v_8_2_2(({n_h_in_acc_psp_lpi_1_dfm
      , conf_info_crt_lpi_1_dfm_160}), (conf_info_rsci_idat_mxwt[23:16]), and_223_cse);
  assign PADDING_LOOP_for_for_index_in_mux_13_nl = MUX_v_16_2_2(({3'b000 , (z_out_1[12:0])}),
      z_out, and_223_cse);
  assign nl_z_out_2 = PADDING_LOOP_for_for_index_in_mux_12_nl * PADDING_LOOP_for_for_index_in_mux_13_nl;
  assign z_out_2 = nl_z_out_2[15:0];

  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [15:0] signext_16_1;
    input [0:0] vector;
  begin
    signext_16_1= {{15{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input [0:0] vector;
  begin
    signext_5_1= {{4{vector[0]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_9_17 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_17 = {{8{vector[8]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_s2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2s_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2s_32_33 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_5_13 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_13 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_16 = vector;
  end
  endfunction


  function automatic [23:0] conv_u2u_24_24 ;
    input [23:0]  vector ;
  begin
    conv_u2u_24_24 = vector;
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute_core
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_inputs_rsc_req_vz,
      plm_inputs_rsc_rls_lz, plm_filters_rsc_req_vz, plm_filters_rsc_rls_lz, plm_outputs_rsc_req_vz,
      plm_outputs_rsc_rls_lz, done_rsc_rdy, done_rsc_vld, plm_inputs_rsci_q_d, plm_inputs_rsci_radr_d,
      plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d, plm_filters_rsci_q_d, plm_filters_rsci_radr_d,
      plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d, plm_outputs_rsci_d_d, plm_outputs_rsci_wadr_d,
      plm_outputs_rsci_we_d_pff
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input plm_inputs_rsc_req_vz;
  output plm_inputs_rsc_rls_lz;
  input plm_filters_rsc_req_vz;
  output plm_filters_rsc_rls_lz;
  input plm_outputs_rsc_req_vz;
  output plm_outputs_rsc_rls_lz;
  input done_rsc_rdy;
  output done_rsc_vld;
  input [31:0] plm_inputs_rsci_q_d;
  output [13:0] plm_inputs_rsci_radr_d;
  output plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] plm_filters_rsci_q_d;
  output [15:0] plm_filters_rsci_radr_d;
  output plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output [31:0] plm_outputs_rsci_d_d;
  output [13:0] plm_outputs_rsci_wadr_d;
  output plm_outputs_rsci_we_d_pff;


  // Interconnect Declarations
  wire core_wen;
  wire conf_info_rsci_bawt;
  wire core_wten;
  wire conf_info_rsci_wen_comp;
  wire [63:0] conf_info_rsci_idat_mxwt;
  wire plm_inputs_rsci_bawt;
  wire [31:0] plm_inputs_rsci_q_d_mxwt;
  wire plm_filters_rsci_bawt;
  wire [31:0] plm_filters_rsci_q_d_mxwt;
  wire plm_outputs_rsci_bawt;
  wire done_rsci_bawt;
  wire done_rsci_wen_comp;
  wire plm_outputs_rsc_rls_obj_bawt;
  wire plm_inputs_rsc_rls_obj_bawt;
  wire plm_filters_rsc_rls_obj_bawt;
  wire plm_filters_rsc_req_obj_bawt;
  reg plm_filters_rsc_req_obj_iswt0;
  wire plm_filters_rsc_req_obj_wen_comp;
  wire plm_inputs_rsc_req_obj_bawt;
  reg plm_inputs_rsc_req_obj_iswt0;
  wire plm_inputs_rsc_req_obj_wen_comp;
  wire plm_outputs_rsc_req_obj_bawt;
  reg plm_outputs_rsc_req_obj_iswt0;
  wire plm_outputs_rsc_req_obj_wen_comp;
  reg CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3;
  reg [29:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4;
  reg CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5;
  wire [1:0] fsm_output;
  wire [4:0] COMPUTE_LOOP_acc_tmp;
  wire [5:0] nl_COMPUTE_LOOP_acc_tmp;
  wire COMPUTE_LOOP_if_COMPUTE_LOOP_if_nand_tmp;
  wire [8:0] operator_8_false_8_acc_tmp;
  wire [9:0] nl_operator_8_false_8_acc_tmp;
  wire [5:0] CONVOLUTION_LOOP_acc_tmp;
  wire [6:0] nl_CONVOLUTION_LOOP_acc_tmp;
  wire CONVOLUTION_LOOP_if_CONVOLUTION_LOOP_if_nand_tmp;
  wire [8:0] operator_8_false_7_acc_tmp;
  wire [9:0] nl_operator_8_false_7_acc_tmp;
  wire [5:0] CONVOLUTION_LOOP_for_acc_tmp;
  wire [6:0] nl_CONVOLUTION_LOOP_for_acc_tmp;
  wire CONVOLUTION_LOOP_for_if_equal_tmp;
  wire [8:0] operator_8_false_5_acc_tmp;
  wire [9:0] nl_operator_8_false_5_acc_tmp;
  wire [8:0] operator_8_false_4_acc_tmp;
  wire [9:0] nl_operator_8_false_4_acc_tmp;
  wire [8:0] operator_8_false_3_acc_tmp;
  wire [9:0] nl_operator_8_false_3_acc_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp;
  wire CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp;
  wire [8:0] operator_8_false_1_acc_tmp;
  wire [9:0] nl_operator_8_false_1_acc_tmp;
  wire COMPUTE_LOOP_COMPUTE_LOOP_or_tmp;
  wire and_9_tmp;
  wire and_7_tmp;
  wire and_5_tmp;
  wire mux_tmp_17;
  wire not_tmp_22;
  wire or_tmp_46;
  wire nand_tmp_7;
  wire mux_tmp_21;
  wire and_dcpl_7;
  wire and_dcpl_11;
  wire and_dcpl_17;
  wire and_dcpl_19;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_32;
  wire and_dcpl_36;
  wire or_dcpl_22;
  wire or_dcpl_31;
  wire and_dcpl_57;
  wire or_dcpl_34;
  wire and_dcpl_59;
  wire or_dcpl_39;
  wire or_dcpl_40;
  wire and_dcpl_66;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_84;
  wire or_tmp_98;
  wire or_tmp_108;
  wire or_tmp_109;
  wire or_tmp_111;
  wire and_113_cse;
  wire exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0;
  wire [3:0] COMPUTE_LOOP_b_4_0_lpi_1_dfm_3_0_1;
  wire exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3_mx0w0;
  wire [4:0] CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_4_0_1;
  wire exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3_mx0w0;
  wire exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0;
  wire [4:0] CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_mx0w0;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6;
  wire exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0;
  reg exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2;
  wire lfst_exit_CONVOLUTION_LOOP_for_for_1_lpi_1_dfm_1;
  reg exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3;
  wire lfst_exit_CONVOLUTION_LOOP_for_1_lpi_1_dfm_1;
  reg exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3;
  reg [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_4_0;
  wire unequal_tmp_1;
  reg exitL_exit_COMPUTE_LOOP_sva;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_1;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_3;
  wire [10:0] COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_3;
  wire CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1;
  reg CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1;
  reg CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0;
  reg [10:0] CONVOLUTION_LOOP_for_for_for_else_mux_itm_1;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1;
  wire CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0;
  wire [44:0] CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0;
  wire CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0;
  wire [48:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1;
  wire [49:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1;
  wire [63:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_9_sdt_sva_1;
  reg exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_3;
  reg main_stage_v_3;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_3;
  reg exit_COMPUTE_LOOP_lpi_1_dfm_2_st_4;
  reg main_stage_v_4;
  reg [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_4;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_2;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2;
  reg [4:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1;
  reg exit_COMPUTE_LOOP_lpi_1_dfm_2;
  reg COMPUTE_LOOP_asn_itm;
  reg exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_1;
  reg exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_2;
  reg exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1;
  reg exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_2;
  reg exit_COMPUTE_LOOP_lpi_1_dfm_2_st_3;
  wire exit_COMPUTE_LOOP_sva_2_mx0w0;
  reg exit_COMPUTE_LOOP_sva_2;
  reg exit_CONVOLUTION_LOOP_lpi_1_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1;
  wire exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0;
  reg exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1;
  wire [48:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1;
  wire [49:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1;
  wire [44:0] CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_45_1_1;
  wire [57:0] CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1;
  wire [58:0] nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1;
  wire [10:0] CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_56_46_1;
  wire and_91_m1c;
  wire and_89_m1c;
  reg reg_conf_info_rsci_iswt0_cse;
  reg reg_plm_filters_rsc_rls_obj_ld_core_psct_cse;
  reg reg_plm_filters_rsc_rls_obj_oswt_cse;
  reg reg_done_rsci_ivld_core_psct_cse;
  reg reg_plm_outputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse;
  reg reg_plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_cse;
  wire COMPUTE_LOOP_buf_acc_data_and_cse;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_6_cse;
  wire COMPUTE_LOOP_and_cse;
  wire CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_2_CONVOLUTION_LOOP_for_for_for_if_2_nor_cse;
  wire nor_55_cse;
  wire nor_40_cse;
  wire and_235_cse;
  wire and_11_cse;
  wire and_10_cse;
  wire or_73_cse;
  wire and_131_cse;
  wire or_113_cse;
  wire CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_if_CONVOLUTION_LOOP_for_if_nor_cse;
  wire CONVOLUTION_LOOP_for_for_if_or_cse;
  wire mux_35_cse;
  reg [13:0] plm_inputs_rsci_radr_d_reg;
  wire [13:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff;
  wire plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  reg [15:0] plm_filters_rsci_radr_d_reg;
  wire [15:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff;
  wire plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff;
  wire [29:0] CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff;
  wire CONVOLUTION_LOOP_for_for_for_if_1_mux_rmff;
  reg [13:0] plm_outputs_rsci_wadr_d_reg;
  wire [13:0] CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff;
  wire plm_outputs_rsci_we_d_iff;
  wire and_50_rmff;
  wire and_34_rmff;
  wire [54:0] CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_5;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_3;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2;
  wire [3:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2;
  wire [7:0] z_out;
  wire [8:0] nl_z_out;
  reg lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1;
  reg [7:0] n_w_out_lpi_1_dfm_1;
  reg [7:0] n_h_out_lpi_1_dfm_1;
  reg [6:0] n_w_in_acc_psp_lpi_1_dfm;
  reg [6:0] n_h_in_acc_psp_lpi_1_dfm;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_1_dfm;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1;
  reg CONVOLUTION_LOOP_for_for_for_acc_0_sva_1;
  reg CONVOLUTION_LOOP_for_for_for_acc_46_sva_1;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_1;
  reg [7:0] CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_1;
  reg [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_2;
  reg [10:0] COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_2;
  reg [44:0] COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_2;
  reg COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_2;
  reg [4:0] CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_4;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm;
  reg exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1;
  reg [15:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1;
  wire [16:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1;
  reg [13:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1;
  wire [14:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1;
  reg [44:0] CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1;
  reg CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1;
  reg [13:0] CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1;
  wire [14:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1;
  reg [13:0] CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2;
  reg CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1;
  reg exit_COMPUTE_LOOP_lpi_1_dfm_2_st_2;
  reg [3:0] COMPUTE_LOOP_b_4_0_lpi_1_3_0;
  reg [7:0] conf_info_crt_lpi_1_dfm_231_224;
  reg conf_info_crt_lpi_1_dfm_192;
  reg conf_info_crt_lpi_1_dfm_160;
  reg [7:0] conf_info_crt_lpi_1_dfm_135_128;
  reg [7:0] conf_info_crt_lpi_1_dfm_103_96;
  reg [7:0] conf_info_crt_lpi_1_dfm_71_64;
  reg [7:0] conf_info_crt_lpi_1_dfm_7_0;
  reg [4:0] CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_2_4_0;
  reg CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1_0;
  wire plm_outputs_rsc_req_obj_iswt0_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire main_stage_v_4_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0;
  wire main_stage_v_1_mx0c1;
  wire [4:0] CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0;
  wire [7:0] conf_info_crt_lpi_1_dfm_231_224_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_71_64_mx0;
  wire [7:0] n_w_out_lpi_1_dfm_3;
  wire [7:0] n_h_out_lpi_1_dfm_3;
  wire [7:0] conf_info_crt_lpi_1_dfm_135_128_mx0;
  wire exit_COMPUTE_LOOP_lpi_1_dfm_2_mx0w0;
  wire [7:0] conf_info_crt_lpi_1_dfm_103_96_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_7_0_mx0;
  wire exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
  wire [6:0] n_w_in_acc_psp_lpi_1_dfm_mx0;
  wire conf_info_crt_lpi_1_dfm_192_mx0;
  wire [6:0] n_h_in_acc_psp_lpi_1_dfm_mx0;
  wire conf_info_crt_lpi_1_dfm_160_mx0;
  wire CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1;
  wire CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1;
  wire COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_1_mx0;
  wire COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_1_mx0;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_3;
  wire [44:0] COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_3;
  wire CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1;
  wire [7:0] if_acc_4_cse_1;
  wire [8:0] nl_if_acc_4_cse_1;
  wire [7:0] pad_sva_1;
  wire signed [16:0] nl_pad_sva_1;
  wire [10:0] else_acc_2_psp_sva_1;
  wire [11:0] nl_else_acc_2_psp_sva_1;
  wire [9:0] else_acc_4_cse_1;
  wire [10:0] nl_else_acc_4_cse_1;
  wire [10:0] else_acc_psp_sva_1;
  wire [11:0] nl_else_acc_psp_sva_1;
  wire [16:0] pad_acc_psp_sva_1;
  wire [17:0] nl_pad_acc_psp_sva_1;
  wire [4:0] CONVOLUTION_LOOP_for_for_i_4_0_sva_2;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2;
  wire [4:0] CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2;
  wire [5:0] nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2;
  wire [3:0] nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2;
  wire [2:0] CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_4;
  wire or_12_cse_1;
  wire or_13_cse_1;
  wire or_4_cse_1;
  wire or_5_cse_1;
  wire or_6_cse_1;
  wire or_7_cse_1;
  wire or_8_cse_1;
  wire or_1_cse_1;
  wire or_2_cse_1;
  wire or_cse_1;
  wire nand_26_cse_1;
  wire nand_15_cse_1;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_mx0;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0;
  wire [7:0] CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1;
  wire [12:0] nl_CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1;
  wire CONVOLUTION_LOOP_for_for_for_asn_3575;
  wire CONVOLUTION_LOOP_for_for_for_asn_3577;
  wire CONVOLUTION_LOOP_for_for_for_asn_3579;
  wire CONVOLUTION_LOOP_for_for_for_asn_3581;
  wire CONVOLUTION_LOOP_for_for_for_asn_3583;
  wire CONVOLUTION_LOOP_for_for_for_asn_3585;
  wire CONVOLUTION_LOOP_for_for_for_asn_3587;
  wire CONVOLUTION_LOOP_for_for_for_asn_3589;
  wire CONVOLUTION_LOOP_for_for_for_asn_3591;
  wire CONVOLUTION_LOOP_for_for_for_asn_3593;
  wire CONVOLUTION_LOOP_for_for_for_asn_3595;
  wire CONVOLUTION_LOOP_for_for_for_asn_3597;
  wire CONVOLUTION_LOOP_for_for_for_asn_3599;
  wire CONVOLUTION_LOOP_for_for_for_asn_3601;
  wire CONVOLUTION_LOOP_for_for_for_asn_3603;
  wire CONVOLUTION_LOOP_for_for_for_asn_3605;
  wire CONVOLUTION_LOOP_for_for_for_asn_3607;
  wire CONVOLUTION_LOOP_for_for_for_asn_3609;
  wire CONVOLUTION_LOOP_for_for_for_asn_3611;
  wire CONVOLUTION_LOOP_for_for_for_asn_3613;
  wire CONVOLUTION_LOOP_for_for_for_asn_3615;
  wire CONVOLUTION_LOOP_for_for_for_asn_3617;
  wire CONVOLUTION_LOOP_for_for_for_asn_3619;
  wire CONVOLUTION_LOOP_for_for_for_asn_3621;
  wire CONVOLUTION_LOOP_for_for_for_asn_3623;
  wire CONVOLUTION_LOOP_for_for_for_asn_3625;
  wire CONVOLUTION_LOOP_for_for_for_asn_3627;
  wire CONVOLUTION_LOOP_for_for_for_asn_3629;
  wire CONVOLUTION_LOOP_for_for_for_asn_3631;
  wire CONVOLUTION_LOOP_for_for_for_asn_3633;
  wire CONVOLUTION_LOOP_for_for_for_asn_3635;
  wire CONVOLUTION_LOOP_for_for_for_asn_3637;
  wire CONVOLUTION_LOOP_for_for_for_asn_3639;
  wire CONVOLUTION_LOOP_for_for_for_asn_3641;
  wire CONVOLUTION_LOOP_for_for_for_asn_3643;
  wire CONVOLUTION_LOOP_for_for_for_asn_3645;
  wire CONVOLUTION_LOOP_for_for_for_asn_3647;
  wire CONVOLUTION_LOOP_for_for_for_asn_3649;
  wire CONVOLUTION_LOOP_for_for_for_asn_3651;
  wire CONVOLUTION_LOOP_for_for_for_asn_3653;
  wire CONVOLUTION_LOOP_for_for_for_asn_3655;
  wire CONVOLUTION_LOOP_for_for_for_asn_3657;
  wire CONVOLUTION_LOOP_for_for_for_asn_3659;
  wire CONVOLUTION_LOOP_for_for_for_asn_3661;
  wire CONVOLUTION_LOOP_for_for_for_asn_3663;
  wire CONVOLUTION_LOOP_for_for_for_asn_3665;
  wire CONVOLUTION_LOOP_for_for_for_asn_3667;
  wire CONVOLUTION_LOOP_for_for_for_asn_3669;
  wire CONVOLUTION_LOOP_for_for_for_asn_3671;
  wire CONVOLUTION_LOOP_for_for_for_asn_3673;
  wire CONVOLUTION_LOOP_for_for_for_asn_3675;
  wire CONVOLUTION_LOOP_for_for_for_asn_3677;
  wire CONVOLUTION_LOOP_for_for_for_asn_3679;
  wire CONVOLUTION_LOOP_for_for_for_asn_3681;
  wire CONVOLUTION_LOOP_for_for_for_asn_3683;
  wire CONVOLUTION_LOOP_for_for_for_asn_3685;
  wire CONVOLUTION_LOOP_for_for_for_asn_3687;
  wire CONVOLUTION_LOOP_for_for_for_asn_3689;
  wire CONVOLUTION_LOOP_for_for_for_asn_3691;
  wire CONVOLUTION_LOOP_for_for_for_asn_3693;
  wire CONVOLUTION_LOOP_for_for_for_asn_3695;
  wire CONVOLUTION_LOOP_for_for_for_asn_3697;
  wire CONVOLUTION_LOOP_for_for_for_asn_3699;
  wire CONVOLUTION_LOOP_for_for_for_asn_3701;
  wire CONVOLUTION_LOOP_for_for_for_asn_3703;
  wire CONVOLUTION_LOOP_for_for_for_asn_3705;
  wire CONVOLUTION_LOOP_for_for_for_asn_3707;
  wire CONVOLUTION_LOOP_for_for_for_asn_3709;
  wire CONVOLUTION_LOOP_for_for_for_asn_3711;
  wire CONVOLUTION_LOOP_for_for_for_asn_3713;
  wire CONVOLUTION_LOOP_for_for_for_asn_3715;
  wire CONVOLUTION_LOOP_for_for_for_asn_3717;
  wire CONVOLUTION_LOOP_for_for_for_asn_3719;
  wire CONVOLUTION_LOOP_for_for_for_asn_3721;
  wire CONVOLUTION_LOOP_for_for_for_asn_3723;
  wire CONVOLUTION_LOOP_for_for_for_asn_3725;
  wire CONVOLUTION_LOOP_for_for_for_asn_3727;
  wire CONVOLUTION_LOOP_for_for_for_asn_3729;
  wire CONVOLUTION_LOOP_for_for_for_asn_3731;
  wire CONVOLUTION_LOOP_for_for_for_asn_3733;
  wire CONVOLUTION_LOOP_for_for_for_asn_3735;
  wire CONVOLUTION_LOOP_for_for_for_asn_3737;
  wire CONVOLUTION_LOOP_for_for_for_asn_3739;
  wire CONVOLUTION_LOOP_for_for_for_asn_3741;
  wire CONVOLUTION_LOOP_for_for_for_asn_3743;
  wire CONVOLUTION_LOOP_for_for_for_asn_3745;
  wire CONVOLUTION_LOOP_for_for_for_asn_3747;
  wire CONVOLUTION_LOOP_for_for_for_asn_3749;
  wire CONVOLUTION_LOOP_for_for_for_asn_3751;
  wire CONVOLUTION_LOOP_for_for_for_asn_3753;
  wire CONVOLUTION_LOOP_for_for_for_asn_3755;
  wire CONVOLUTION_LOOP_for_for_for_asn_3757;
  wire CONVOLUTION_LOOP_for_for_for_asn_3759;
  wire CONVOLUTION_LOOP_for_for_for_asn_3761;
  wire CONVOLUTION_LOOP_for_for_for_asn_3763;
  wire CONVOLUTION_LOOP_for_for_for_asn_3765;
  wire CONVOLUTION_LOOP_for_for_for_asn_3767;
  wire CONVOLUTION_LOOP_for_for_for_asn_3769;
  wire CONVOLUTION_LOOP_for_for_for_asn_3771;
  wire CONVOLUTION_LOOP_for_for_for_asn_3773;
  wire CONVOLUTION_LOOP_for_for_for_asn_3775;
  wire CONVOLUTION_LOOP_for_for_for_asn_3777;
  wire CONVOLUTION_LOOP_for_for_for_asn_3779;
  wire CONVOLUTION_LOOP_for_for_for_asn_3781;
  wire CONVOLUTION_LOOP_for_for_for_asn_3783;
  wire CONVOLUTION_LOOP_for_for_for_asn_3785;
  wire CONVOLUTION_LOOP_for_for_for_asn_3787;
  wire CONVOLUTION_LOOP_for_for_for_asn_3789;
  wire CONVOLUTION_LOOP_for_for_for_asn_3791;
  wire CONVOLUTION_LOOP_for_for_for_asn_3793;
  wire CONVOLUTION_LOOP_for_for_for_asn_3795;
  wire CONVOLUTION_LOOP_for_for_for_asn_3797;
  wire CONVOLUTION_LOOP_for_for_for_asn_3799;
  wire CONVOLUTION_LOOP_for_for_for_asn_3801;
  wire CONVOLUTION_LOOP_for_for_for_asn_3803;
  wire CONVOLUTION_LOOP_for_for_for_asn_3805;
  wire CONVOLUTION_LOOP_for_for_for_asn_3807;
  wire CONVOLUTION_LOOP_for_for_for_asn_3809;
  wire CONVOLUTION_LOOP_for_for_for_asn_3811;
  wire CONVOLUTION_LOOP_for_for_for_asn_3813;
  wire CONVOLUTION_LOOP_for_for_for_asn_3815;
  wire CONVOLUTION_LOOP_for_for_for_asn_3817;
  wire CONVOLUTION_LOOP_for_for_for_asn_3819;
  wire CONVOLUTION_LOOP_for_for_for_asn_3821;
  wire CONVOLUTION_LOOP_for_for_for_asn_3823;
  wire CONVOLUTION_LOOP_for_for_for_asn_3825;
  wire CONVOLUTION_LOOP_for_for_for_asn_3827;
  wire CONVOLUTION_LOOP_for_for_for_asn_3829;
  wire CONVOLUTION_LOOP_for_for_for_asn_3831;
  wire CONVOLUTION_LOOP_for_for_for_asn_3833;
  wire CONVOLUTION_LOOP_for_for_for_asn_3835;
  wire CONVOLUTION_LOOP_for_for_for_asn_3837;
  wire CONVOLUTION_LOOP_for_for_for_asn_3839;
  wire CONVOLUTION_LOOP_for_for_for_asn_3841;
  wire CONVOLUTION_LOOP_for_for_for_asn_3843;
  wire CONVOLUTION_LOOP_for_for_for_asn_3845;
  wire CONVOLUTION_LOOP_for_for_for_asn_3847;
  wire CONVOLUTION_LOOP_for_for_for_asn_3849;
  wire CONVOLUTION_LOOP_for_for_for_asn_3851;
  wire CONVOLUTION_LOOP_for_for_for_asn_3853;
  wire CONVOLUTION_LOOP_for_for_for_asn_3855;
  wire CONVOLUTION_LOOP_for_for_for_asn_3857;
  wire CONVOLUTION_LOOP_for_for_for_asn_3859;
  wire CONVOLUTION_LOOP_for_for_for_asn_3861;
  wire CONVOLUTION_LOOP_for_for_for_asn_3863;
  wire CONVOLUTION_LOOP_for_for_for_asn_3865;
  wire CONVOLUTION_LOOP_for_for_for_asn_3867;
  wire CONVOLUTION_LOOP_for_for_for_asn_3869;
  wire CONVOLUTION_LOOP_for_for_for_asn_3871;
  wire CONVOLUTION_LOOP_for_for_for_asn_3873;
  wire CONVOLUTION_LOOP_for_for_for_asn_3875;
  wire CONVOLUTION_LOOP_for_for_for_asn_3877;
  wire CONVOLUTION_LOOP_for_for_for_asn_3879;
  wire CONVOLUTION_LOOP_for_for_for_asn_3881;
  wire CONVOLUTION_LOOP_for_for_for_asn_3883;
  wire CONVOLUTION_LOOP_for_for_for_asn_3885;
  wire CONVOLUTION_LOOP_for_for_for_asn_3887;
  wire CONVOLUTION_LOOP_for_for_for_asn_3889;
  wire CONVOLUTION_LOOP_for_for_for_asn_3891;
  wire CONVOLUTION_LOOP_for_for_for_asn_3893;
  wire CONVOLUTION_LOOP_for_for_for_asn_3895;
  wire CONVOLUTION_LOOP_for_for_for_asn_3897;
  wire CONVOLUTION_LOOP_for_for_for_asn_3899;
  wire CONVOLUTION_LOOP_for_for_for_asn_3901;
  wire CONVOLUTION_LOOP_for_for_for_asn_3903;
  wire CONVOLUTION_LOOP_for_for_for_asn_3905;
  wire CONVOLUTION_LOOP_for_for_for_asn_3907;
  wire CONVOLUTION_LOOP_for_for_for_asn_3909;
  wire CONVOLUTION_LOOP_for_for_for_asn_3911;
  wire CONVOLUTION_LOOP_for_for_for_asn_3913;
  wire CONVOLUTION_LOOP_for_for_for_asn_3915;
  wire CONVOLUTION_LOOP_for_for_for_asn_3917;
  wire CONVOLUTION_LOOP_for_for_for_asn_3919;
  wire CONVOLUTION_LOOP_for_for_for_asn_3921;
  wire CONVOLUTION_LOOP_for_for_for_asn_3923;
  wire CONVOLUTION_LOOP_for_for_for_asn_3925;
  wire CONVOLUTION_LOOP_for_for_for_asn_3927;
  wire CONVOLUTION_LOOP_for_for_for_asn_3929;
  wire CONVOLUTION_LOOP_for_for_for_asn_3931;
  wire CONVOLUTION_LOOP_for_for_for_asn_3933;
  wire CONVOLUTION_LOOP_for_for_for_asn_3935;
  wire CONVOLUTION_LOOP_for_for_for_asn_3937;
  wire CONVOLUTION_LOOP_for_for_for_asn_3939;
  wire CONVOLUTION_LOOP_for_for_for_asn_3941;
  wire CONVOLUTION_LOOP_for_for_for_asn_3943;
  wire CONVOLUTION_LOOP_for_for_for_asn_3945;
  wire CONVOLUTION_LOOP_for_for_for_asn_3947;
  wire CONVOLUTION_LOOP_for_for_for_asn_3949;
  wire CONVOLUTION_LOOP_for_for_for_asn_3951;
  wire CONVOLUTION_LOOP_for_for_for_asn_3953;
  wire CONVOLUTION_LOOP_for_for_for_asn_3955;
  wire CONVOLUTION_LOOP_for_for_for_asn_3957;
  wire CONVOLUTION_LOOP_for_for_for_asn_3959;
  wire CONVOLUTION_LOOP_for_for_for_asn_3961;
  wire CONVOLUTION_LOOP_for_for_for_asn_3963;
  wire CONVOLUTION_LOOP_for_for_for_asn_3965;
  wire CONVOLUTION_LOOP_for_for_for_asn_3967;
  wire CONVOLUTION_LOOP_for_for_for_asn_3969;
  wire CONVOLUTION_LOOP_for_for_for_asn_3971;
  wire CONVOLUTION_LOOP_for_for_for_asn_3973;
  wire CONVOLUTION_LOOP_for_for_for_asn_3975;
  wire CONVOLUTION_LOOP_for_for_for_asn_3977;
  wire CONVOLUTION_LOOP_for_for_for_asn_3979;
  wire CONVOLUTION_LOOP_for_for_for_asn_3981;
  wire CONVOLUTION_LOOP_for_for_for_asn_3983;
  wire CONVOLUTION_LOOP_for_for_for_asn_3985;
  wire CONVOLUTION_LOOP_for_for_for_asn_3987;
  wire CONVOLUTION_LOOP_for_for_for_asn_3989;
  wire CONVOLUTION_LOOP_for_for_for_asn_3991;
  wire CONVOLUTION_LOOP_for_for_for_asn_3993;
  wire CONVOLUTION_LOOP_for_for_for_asn_3995;
  wire CONVOLUTION_LOOP_for_for_for_asn_3997;
  wire CONVOLUTION_LOOP_for_for_for_asn_3999;
  wire CONVOLUTION_LOOP_for_for_for_asn_4001;
  wire CONVOLUTION_LOOP_for_for_for_asn_4003;
  wire CONVOLUTION_LOOP_for_for_for_asn_4005;
  wire CONVOLUTION_LOOP_for_for_for_asn_4007;
  wire CONVOLUTION_LOOP_for_for_for_asn_4009;
  wire CONVOLUTION_LOOP_for_for_for_asn_4011;
  wire CONVOLUTION_LOOP_for_for_for_asn_4013;
  wire CONVOLUTION_LOOP_for_for_for_asn_4015;
  wire CONVOLUTION_LOOP_for_for_for_asn_4017;
  wire CONVOLUTION_LOOP_for_for_for_asn_4019;
  wire CONVOLUTION_LOOP_for_for_for_asn_4021;
  wire CONVOLUTION_LOOP_for_for_for_asn_4023;
  wire CONVOLUTION_LOOP_for_for_for_asn_4025;
  wire CONVOLUTION_LOOP_for_for_for_asn_4027;
  wire CONVOLUTION_LOOP_for_for_for_asn_4029;
  wire CONVOLUTION_LOOP_for_for_for_asn_4031;
  wire CONVOLUTION_LOOP_for_for_for_asn_4033;
  wire CONVOLUTION_LOOP_for_for_for_asn_4035;
  wire CONVOLUTION_LOOP_for_for_for_asn_4037;
  wire CONVOLUTION_LOOP_for_for_for_asn_4039;
  wire CONVOLUTION_LOOP_for_for_for_asn_4041;
  wire CONVOLUTION_LOOP_for_for_for_asn_4043;
  wire CONVOLUTION_LOOP_for_for_for_asn_4045;
  wire CONVOLUTION_LOOP_for_for_for_asn_4047;
  wire CONVOLUTION_LOOP_for_for_for_asn_4049;
  wire CONVOLUTION_LOOP_for_for_for_asn_4051;
  wire CONVOLUTION_LOOP_for_for_for_asn_4053;
  wire CONVOLUTION_LOOP_for_for_for_asn_4055;
  wire CONVOLUTION_LOOP_for_for_for_asn_4057;
  wire CONVOLUTION_LOOP_for_for_for_asn_4059;
  wire CONVOLUTION_LOOP_for_for_for_asn_4061;
  wire CONVOLUTION_LOOP_for_for_for_asn_4063;
  wire CONVOLUTION_LOOP_for_for_for_asn_4065;
  wire CONVOLUTION_LOOP_for_for_for_asn_4067;
  wire CONVOLUTION_LOOP_for_for_for_asn_4069;
  wire CONVOLUTION_LOOP_for_for_for_asn_4071;
  wire CONVOLUTION_LOOP_for_for_for_asn_4073;
  wire CONVOLUTION_LOOP_for_for_for_asn_4075;
  wire CONVOLUTION_LOOP_for_for_for_asn_4077;
  wire CONVOLUTION_LOOP_for_for_for_asn_4079;
  wire CONVOLUTION_LOOP_for_for_for_asn_4081;
  wire CONVOLUTION_LOOP_for_for_for_asn_4083;
  wire CONVOLUTION_LOOP_for_for_for_asn_4085;
  wire CONVOLUTION_LOOP_for_for_for_asn_4087;
  wire CONVOLUTION_LOOP_for_for_for_asn_4089;
  wire CONVOLUTION_LOOP_for_for_for_asn_4091;
  wire CONVOLUTION_LOOP_for_for_for_asn_4093;
  wire CONVOLUTION_LOOP_for_for_for_asn_4095;
  wire CONVOLUTION_LOOP_for_for_for_asn_4097;
  wire CONVOLUTION_LOOP_for_for_for_asn_4099;
  wire CONVOLUTION_LOOP_for_for_for_asn_4101;
  wire CONVOLUTION_LOOP_for_for_for_asn_4103;
  wire CONVOLUTION_LOOP_for_for_for_asn_4105;
  wire CONVOLUTION_LOOP_for_for_for_asn_4107;
  wire CONVOLUTION_LOOP_for_for_for_asn_4109;
  wire CONVOLUTION_LOOP_for_for_for_asn_4111;
  wire CONVOLUTION_LOOP_for_for_for_asn_4113;
  wire CONVOLUTION_LOOP_for_for_for_asn_4115;
  wire CONVOLUTION_LOOP_for_for_for_asn_4117;
  wire CONVOLUTION_LOOP_for_for_for_asn_4119;
  wire CONVOLUTION_LOOP_for_for_for_asn_4121;
  wire CONVOLUTION_LOOP_for_for_for_asn_4123;
  wire CONVOLUTION_LOOP_for_for_for_asn_4125;
  wire CONVOLUTION_LOOP_for_for_for_asn_4127;
  wire CONVOLUTION_LOOP_for_for_for_asn_4129;
  wire CONVOLUTION_LOOP_for_for_for_asn_4131;
  wire CONVOLUTION_LOOP_for_for_for_asn_4133;
  wire CONVOLUTION_LOOP_for_for_for_asn_4135;
  wire CONVOLUTION_LOOP_for_for_for_asn_4137;
  wire CONVOLUTION_LOOP_for_for_for_asn_4139;
  wire CONVOLUTION_LOOP_for_for_for_asn_4141;
  wire CONVOLUTION_LOOP_for_for_for_asn_4143;
  wire CONVOLUTION_LOOP_for_for_for_asn_4145;
  wire CONVOLUTION_LOOP_for_for_for_asn_4147;
  wire CONVOLUTION_LOOP_for_for_for_asn_4149;
  wire CONVOLUTION_LOOP_for_for_for_asn_4151;
  wire CONVOLUTION_LOOP_for_for_for_asn_4153;
  wire CONVOLUTION_LOOP_for_for_for_asn_4155;
  wire CONVOLUTION_LOOP_for_for_for_asn_4157;
  wire CONVOLUTION_LOOP_for_for_for_asn_4159;
  wire CONVOLUTION_LOOP_for_for_for_asn_4161;
  wire CONVOLUTION_LOOP_for_for_for_asn_4163;
  wire CONVOLUTION_LOOP_for_for_for_asn_4165;
  wire CONVOLUTION_LOOP_for_for_for_asn_4167;
  wire CONVOLUTION_LOOP_for_for_for_asn_4169;
  wire CONVOLUTION_LOOP_for_for_for_asn_4171;
  wire CONVOLUTION_LOOP_for_for_for_asn_4173;
  wire CONVOLUTION_LOOP_for_for_for_asn_4175;
  wire CONVOLUTION_LOOP_for_for_for_asn_4177;
  wire CONVOLUTION_LOOP_for_for_for_asn_4179;
  wire CONVOLUTION_LOOP_for_for_for_asn_4181;
  wire CONVOLUTION_LOOP_for_for_for_asn_4183;
  wire CONVOLUTION_LOOP_for_for_for_asn_4185;
  wire CONVOLUTION_LOOP_for_for_for_asn_4187;
  wire CONVOLUTION_LOOP_for_for_for_asn_4189;
  wire CONVOLUTION_LOOP_for_for_for_asn_4191;
  wire CONVOLUTION_LOOP_for_for_for_asn_4193;
  wire CONVOLUTION_LOOP_for_for_for_asn_4195;
  wire CONVOLUTION_LOOP_for_for_for_asn_4197;
  wire CONVOLUTION_LOOP_for_for_for_asn_4199;
  wire CONVOLUTION_LOOP_for_for_for_asn_4201;
  wire CONVOLUTION_LOOP_for_for_for_asn_4203;
  wire CONVOLUTION_LOOP_for_for_for_asn_4205;
  wire CONVOLUTION_LOOP_for_for_for_asn_4207;
  wire CONVOLUTION_LOOP_for_for_for_asn_4209;
  wire CONVOLUTION_LOOP_for_for_for_asn_4211;
  wire CONVOLUTION_LOOP_for_for_for_asn_4213;
  wire CONVOLUTION_LOOP_for_for_for_asn_4215;
  wire CONVOLUTION_LOOP_for_for_for_asn_4217;
  wire CONVOLUTION_LOOP_for_for_for_asn_4219;
  wire CONVOLUTION_LOOP_for_for_for_asn_4221;
  wire CONVOLUTION_LOOP_for_for_for_asn_4223;
  wire CONVOLUTION_LOOP_for_for_for_asn_4225;
  wire CONVOLUTION_LOOP_for_for_for_asn_4227;
  wire CONVOLUTION_LOOP_for_for_for_asn_4229;
  wire CONVOLUTION_LOOP_for_for_for_asn_4231;
  wire CONVOLUTION_LOOP_for_for_for_asn_4233;
  wire CONVOLUTION_LOOP_for_for_for_asn_4235;
  wire CONVOLUTION_LOOP_for_for_for_asn_4237;
  wire CONVOLUTION_LOOP_for_for_for_asn_4239;
  wire CONVOLUTION_LOOP_for_for_for_asn_4241;
  wire CONVOLUTION_LOOP_for_for_for_asn_4243;
  wire CONVOLUTION_LOOP_for_for_for_asn_4245;
  wire CONVOLUTION_LOOP_for_for_for_asn_4247;
  wire CONVOLUTION_LOOP_for_for_for_asn_4249;
  wire CONVOLUTION_LOOP_for_for_for_asn_4251;
  wire CONVOLUTION_LOOP_for_for_for_asn_4253;
  wire CONVOLUTION_LOOP_for_for_for_asn_4255;
  wire CONVOLUTION_LOOP_for_for_for_asn_4257;
  wire CONVOLUTION_LOOP_for_for_for_asn_4259;
  wire CONVOLUTION_LOOP_for_for_for_asn_4261;
  wire CONVOLUTION_LOOP_for_for_for_asn_4263;
  wire CONVOLUTION_LOOP_for_for_for_asn_4265;
  wire CONVOLUTION_LOOP_for_for_for_asn_4267;
  wire CONVOLUTION_LOOP_for_for_for_asn_4269;
  wire CONVOLUTION_LOOP_for_for_for_asn_4271;
  wire CONVOLUTION_LOOP_for_for_for_asn_4273;
  wire CONVOLUTION_LOOP_for_for_for_asn_4275;
  wire CONVOLUTION_LOOP_for_for_for_asn_4277;
  wire CONVOLUTION_LOOP_for_for_for_asn_4279;
  wire CONVOLUTION_LOOP_for_for_for_asn_4281;
  wire CONVOLUTION_LOOP_for_for_for_asn_4283;
  wire CONVOLUTION_LOOP_for_for_for_asn_4285;
  wire CONVOLUTION_LOOP_for_for_for_asn_4287;
  wire CONVOLUTION_LOOP_for_for_for_asn_4289;
  wire CONVOLUTION_LOOP_for_for_for_asn_4291;
  wire CONVOLUTION_LOOP_for_for_for_asn_4293;
  wire CONVOLUTION_LOOP_for_for_for_asn_4295;
  wire CONVOLUTION_LOOP_for_for_for_asn_4297;
  wire CONVOLUTION_LOOP_for_for_for_asn_4299;
  wire CONVOLUTION_LOOP_for_for_for_asn_4301;
  wire CONVOLUTION_LOOP_for_for_for_asn_4303;
  wire CONVOLUTION_LOOP_for_for_for_asn_4305;
  wire CONVOLUTION_LOOP_for_for_for_asn_4307;
  wire CONVOLUTION_LOOP_for_for_for_asn_4309;
  wire CONVOLUTION_LOOP_for_for_for_asn_4311;
  wire CONVOLUTION_LOOP_for_for_for_asn_4313;
  wire CONVOLUTION_LOOP_for_for_for_asn_4315;
  wire CONVOLUTION_LOOP_for_for_for_asn_4317;
  wire CONVOLUTION_LOOP_for_for_for_asn_4319;
  wire CONVOLUTION_LOOP_for_for_for_asn_4321;
  wire CONVOLUTION_LOOP_for_for_for_asn_4323;
  wire CONVOLUTION_LOOP_for_for_for_asn_4325;
  wire CONVOLUTION_LOOP_for_for_for_asn_4327;
  wire CONVOLUTION_LOOP_for_for_for_asn_4329;
  wire CONVOLUTION_LOOP_for_for_for_asn_4331;
  wire CONVOLUTION_LOOP_for_for_for_asn_4333;
  wire CONVOLUTION_LOOP_for_for_for_asn_4335;
  wire CONVOLUTION_LOOP_for_for_for_asn_4337;
  wire CONVOLUTION_LOOP_for_for_for_asn_4339;
  wire CONVOLUTION_LOOP_for_for_for_asn_4341;
  wire CONVOLUTION_LOOP_for_for_for_asn_4343;
  wire CONVOLUTION_LOOP_for_for_for_asn_4345;
  wire CONVOLUTION_LOOP_for_for_for_asn_4347;
  wire CONVOLUTION_LOOP_for_for_for_asn_4349;
  wire CONVOLUTION_LOOP_for_for_for_asn_4351;
  wire CONVOLUTION_LOOP_for_for_for_asn_4353;
  wire CONVOLUTION_LOOP_for_for_for_asn_4355;
  wire CONVOLUTION_LOOP_for_for_for_asn_4357;
  wire CONVOLUTION_LOOP_for_for_for_asn_4359;
  wire CONVOLUTION_LOOP_for_for_for_asn_4361;
  wire CONVOLUTION_LOOP_for_for_for_asn_4363;
  wire CONVOLUTION_LOOP_for_for_for_asn_4365;
  wire CONVOLUTION_LOOP_for_for_for_asn_4367;
  wire CONVOLUTION_LOOP_for_for_for_asn_4369;
  wire CONVOLUTION_LOOP_for_for_for_asn_4371;
  wire CONVOLUTION_LOOP_for_for_for_asn_4373;
  wire CONVOLUTION_LOOP_for_for_for_asn_4375;
  wire CONVOLUTION_LOOP_for_for_for_asn_4377;
  wire CONVOLUTION_LOOP_for_for_for_asn_4379;
  wire CONVOLUTION_LOOP_for_for_for_asn_4381;
  wire CONVOLUTION_LOOP_for_for_for_asn_4383;
  wire CONVOLUTION_LOOP_for_for_for_asn_4385;
  wire CONVOLUTION_LOOP_for_for_for_asn_4387;
  wire CONVOLUTION_LOOP_for_for_for_asn_4389;
  wire CONVOLUTION_LOOP_for_for_for_asn_4391;
  wire CONVOLUTION_LOOP_for_for_for_asn_4393;
  wire CONVOLUTION_LOOP_for_for_for_asn_4395;
  wire CONVOLUTION_LOOP_for_for_for_asn_4397;
  wire CONVOLUTION_LOOP_for_for_for_asn_4399;
  wire CONVOLUTION_LOOP_for_for_for_asn_4401;
  wire CONVOLUTION_LOOP_for_for_for_asn_4403;
  wire CONVOLUTION_LOOP_for_for_for_asn_4405;
  wire CONVOLUTION_LOOP_for_for_for_asn_4407;
  wire CONVOLUTION_LOOP_for_for_for_asn_4409;
  wire CONVOLUTION_LOOP_for_for_for_asn_4411;
  wire CONVOLUTION_LOOP_for_for_for_asn_4413;
  wire CONVOLUTION_LOOP_for_for_for_asn_4415;
  wire CONVOLUTION_LOOP_for_for_for_asn_4417;
  wire CONVOLUTION_LOOP_for_for_for_asn_4419;
  wire CONVOLUTION_LOOP_for_for_for_asn_4421;
  wire CONVOLUTION_LOOP_for_for_for_asn_4423;
  wire CONVOLUTION_LOOP_for_for_for_asn_4425;
  wire CONVOLUTION_LOOP_for_for_for_asn_4427;
  wire CONVOLUTION_LOOP_for_for_for_asn_4429;
  wire CONVOLUTION_LOOP_for_for_for_asn_4431;
  wire CONVOLUTION_LOOP_for_for_for_asn_4433;
  wire CONVOLUTION_LOOP_for_for_for_asn_4435;
  wire CONVOLUTION_LOOP_for_for_for_asn_4437;
  wire CONVOLUTION_LOOP_for_for_for_asn_4439;
  wire CONVOLUTION_LOOP_for_for_for_asn_4441;
  wire CONVOLUTION_LOOP_for_for_for_asn_4443;
  wire CONVOLUTION_LOOP_for_for_for_asn_4445;
  wire CONVOLUTION_LOOP_for_for_for_asn_4447;
  wire CONVOLUTION_LOOP_for_for_for_asn_4449;
  wire CONVOLUTION_LOOP_for_for_for_asn_4451;
  wire CONVOLUTION_LOOP_for_for_for_asn_4453;
  wire CONVOLUTION_LOOP_for_for_for_asn_4455;
  wire CONVOLUTION_LOOP_for_for_for_asn_4457;
  wire CONVOLUTION_LOOP_for_for_for_asn_4459;
  wire CONVOLUTION_LOOP_for_for_for_asn_4461;
  wire CONVOLUTION_LOOP_for_for_for_asn_4463;
  wire CONVOLUTION_LOOP_for_for_for_asn_4465;
  wire CONVOLUTION_LOOP_for_for_for_asn_4467;
  wire CONVOLUTION_LOOP_for_for_for_asn_4469;
  wire CONVOLUTION_LOOP_for_for_for_asn_4471;
  wire CONVOLUTION_LOOP_for_for_for_asn_4473;
  wire CONVOLUTION_LOOP_for_for_for_asn_4475;
  wire CONVOLUTION_LOOP_for_for_for_asn_4477;
  wire CONVOLUTION_LOOP_for_for_for_asn_4479;
  wire CONVOLUTION_LOOP_for_for_for_asn_4481;
  wire CONVOLUTION_LOOP_for_for_for_asn_4483;
  wire CONVOLUTION_LOOP_for_for_for_asn_4485;
  wire CONVOLUTION_LOOP_for_for_for_asn_4487;
  wire CONVOLUTION_LOOP_for_for_for_asn_4489;
  wire CONVOLUTION_LOOP_for_for_for_asn_4491;
  wire CONVOLUTION_LOOP_for_for_for_asn_4493;
  wire CONVOLUTION_LOOP_for_for_for_asn_4495;
  wire CONVOLUTION_LOOP_for_for_for_asn_4497;
  wire CONVOLUTION_LOOP_for_for_for_asn_4499;
  wire CONVOLUTION_LOOP_for_for_for_asn_4501;
  wire CONVOLUTION_LOOP_for_for_for_asn_4503;
  wire CONVOLUTION_LOOP_for_for_for_asn_4505;
  wire CONVOLUTION_LOOP_for_for_for_asn_4507;
  wire CONVOLUTION_LOOP_for_for_for_asn_4509;
  wire CONVOLUTION_LOOP_for_for_for_asn_4511;
  wire CONVOLUTION_LOOP_for_for_for_asn_4513;
  wire CONVOLUTION_LOOP_for_for_for_asn_4515;
  wire CONVOLUTION_LOOP_for_for_for_asn_4517;
  wire CONVOLUTION_LOOP_for_for_for_asn_4519;
  wire CONVOLUTION_LOOP_for_for_for_asn_4521;
  wire CONVOLUTION_LOOP_for_for_for_asn_4523;
  wire CONVOLUTION_LOOP_for_for_for_asn_4525;
  wire CONVOLUTION_LOOP_for_for_for_asn_4527;
  wire CONVOLUTION_LOOP_for_for_for_asn_4529;
  wire CONVOLUTION_LOOP_for_for_for_asn_4531;
  wire CONVOLUTION_LOOP_for_for_for_asn_4533;
  wire CONVOLUTION_LOOP_for_for_for_asn_4535;
  wire CONVOLUTION_LOOP_for_for_for_asn_4537;
  wire CONVOLUTION_LOOP_for_for_for_asn_4539;
  wire CONVOLUTION_LOOP_for_for_for_asn_4541;
  wire CONVOLUTION_LOOP_for_for_for_asn_4543;
  wire CONVOLUTION_LOOP_for_for_for_asn_4545;
  wire CONVOLUTION_LOOP_for_for_for_asn_4547;
  wire CONVOLUTION_LOOP_for_for_for_asn_4549;
  wire CONVOLUTION_LOOP_for_for_for_asn_4551;
  wire CONVOLUTION_LOOP_for_for_for_asn_4553;
  wire CONVOLUTION_LOOP_for_for_for_asn_4555;
  wire CONVOLUTION_LOOP_for_for_for_asn_4557;
  wire CONVOLUTION_LOOP_for_for_for_asn_4559;
  wire CONVOLUTION_LOOP_for_for_for_asn_4561;
  wire CONVOLUTION_LOOP_for_for_for_asn_4563;
  wire CONVOLUTION_LOOP_for_for_for_asn_4565;
  wire CONVOLUTION_LOOP_for_for_for_asn_4567;
  wire CONVOLUTION_LOOP_for_for_for_asn_4569;
  wire CONVOLUTION_LOOP_for_for_for_asn_4571;
  wire CONVOLUTION_LOOP_for_for_for_asn_4573;
  wire CONVOLUTION_LOOP_for_for_for_asn_4575;
  wire CONVOLUTION_LOOP_for_for_for_asn_4577;
  wire CONVOLUTION_LOOP_for_for_for_asn_4579;
  wire CONVOLUTION_LOOP_for_for_for_asn_4581;
  wire CONVOLUTION_LOOP_for_for_for_asn_4583;
  wire CONVOLUTION_LOOP_for_for_for_asn_4585;
  wire CONVOLUTION_LOOP_for_for_for_asn_4587;
  wire CONVOLUTION_LOOP_for_for_for_asn_4589;
  wire CONVOLUTION_LOOP_for_for_for_asn_4591;
  wire CONVOLUTION_LOOP_for_for_for_asn_4593;
  wire CONVOLUTION_LOOP_for_for_for_asn_4595;
  wire CONVOLUTION_LOOP_for_for_for_asn_4597;
  wire CONVOLUTION_LOOP_for_for_for_asn_4599;
  wire CONVOLUTION_LOOP_for_for_for_asn_4601;
  wire CONVOLUTION_LOOP_for_for_for_asn_4603;
  wire CONVOLUTION_LOOP_for_for_for_asn_4605;
  wire CONVOLUTION_LOOP_for_for_for_asn_4607;
  wire CONVOLUTION_LOOP_for_for_for_asn_4609;
  wire CONVOLUTION_LOOP_for_for_for_asn_4611;
  wire CONVOLUTION_LOOP_for_for_for_asn_4613;
  wire CONVOLUTION_LOOP_for_for_for_asn_4615;
  wire CONVOLUTION_LOOP_for_for_for_asn_4617;
  wire CONVOLUTION_LOOP_for_for_for_asn_4619;
  wire CONVOLUTION_LOOP_for_for_for_asn_4621;
  wire CONVOLUTION_LOOP_for_for_for_asn_4623;
  wire CONVOLUTION_LOOP_for_for_for_asn_4625;
  wire CONVOLUTION_LOOP_for_for_for_asn_4627;
  wire CONVOLUTION_LOOP_for_for_for_asn_4629;
  wire CONVOLUTION_LOOP_for_for_for_asn_4631;
  wire CONVOLUTION_LOOP_for_for_for_asn_4633;
  wire CONVOLUTION_LOOP_for_for_for_asn_4635;
  wire CONVOLUTION_LOOP_for_for_for_asn_4637;
  wire CONVOLUTION_LOOP_for_for_for_asn_4639;
  wire CONVOLUTION_LOOP_for_for_for_asn_4641;
  wire CONVOLUTION_LOOP_for_for_for_asn_4643;
  wire CONVOLUTION_LOOP_for_for_for_asn_4645;
  wire CONVOLUTION_LOOP_for_for_for_asn_4647;
  wire CONVOLUTION_LOOP_for_for_for_asn_4649;
  wire CONVOLUTION_LOOP_for_for_for_asn_4651;
  wire CONVOLUTION_LOOP_for_for_for_asn_4653;
  wire CONVOLUTION_LOOP_for_for_for_asn_4655;
  wire CONVOLUTION_LOOP_for_for_for_asn_4657;
  wire CONVOLUTION_LOOP_for_for_for_asn_4659;
  wire CONVOLUTION_LOOP_for_for_for_asn_4661;
  wire CONVOLUTION_LOOP_for_for_for_asn_4663;
  wire CONVOLUTION_LOOP_for_for_for_asn_4665;
  wire CONVOLUTION_LOOP_for_for_for_asn_4667;
  wire CONVOLUTION_LOOP_for_for_for_asn_4669;
  wire CONVOLUTION_LOOP_for_for_for_asn_4671;
  wire CONVOLUTION_LOOP_for_for_for_asn_4673;
  wire CONVOLUTION_LOOP_for_for_for_asn_4675;
  wire CONVOLUTION_LOOP_for_for_for_asn_4677;
  wire CONVOLUTION_LOOP_for_for_for_asn_4679;
  wire CONVOLUTION_LOOP_for_for_for_asn_4681;
  wire CONVOLUTION_LOOP_for_for_for_asn_4683;
  wire CONVOLUTION_LOOP_for_for_for_asn_4685;
  wire CONVOLUTION_LOOP_for_for_for_asn_4687;
  wire CONVOLUTION_LOOP_for_for_for_asn_4689;
  wire CONVOLUTION_LOOP_for_for_for_asn_4691;
  wire CONVOLUTION_LOOP_for_for_for_asn_4693;
  wire CONVOLUTION_LOOP_for_for_for_asn_4695;
  wire CONVOLUTION_LOOP_for_for_for_asn_4697;
  wire CONVOLUTION_LOOP_for_for_for_asn_4699;
  wire CONVOLUTION_LOOP_for_for_for_asn_4701;
  wire CONVOLUTION_LOOP_for_for_for_asn_4703;
  wire CONVOLUTION_LOOP_for_for_for_asn_4705;
  wire CONVOLUTION_LOOP_for_for_for_asn_4707;
  wire CONVOLUTION_LOOP_for_for_for_asn_4709;
  wire CONVOLUTION_LOOP_for_for_for_asn_4711;
  wire CONVOLUTION_LOOP_for_for_for_asn_4713;
  wire CONVOLUTION_LOOP_for_for_for_asn_4715;
  wire CONVOLUTION_LOOP_for_for_for_asn_4717;
  wire CONVOLUTION_LOOP_for_for_for_asn_4719;
  wire CONVOLUTION_LOOP_for_for_for_asn_4721;
  wire CONVOLUTION_LOOP_for_for_for_asn_4723;
  wire CONVOLUTION_LOOP_for_for_for_asn_4725;
  wire CONVOLUTION_LOOP_for_for_for_asn_4727;
  wire CONVOLUTION_LOOP_for_for_for_asn_4729;
  wire CONVOLUTION_LOOP_for_for_for_asn_4731;
  wire CONVOLUTION_LOOP_for_for_for_asn_4733;
  wire CONVOLUTION_LOOP_for_for_for_asn_4735;
  wire CONVOLUTION_LOOP_for_for_for_asn_4737;
  wire CONVOLUTION_LOOP_for_for_for_asn_4739;
  wire CONVOLUTION_LOOP_for_for_for_asn_4741;
  wire CONVOLUTION_LOOP_for_for_for_asn_4743;
  wire CONVOLUTION_LOOP_for_for_for_asn_4745;
  wire CONVOLUTION_LOOP_for_for_for_asn_4747;
  wire CONVOLUTION_LOOP_for_for_for_asn_4749;
  wire CONVOLUTION_LOOP_for_for_for_asn_4751;
  wire CONVOLUTION_LOOP_for_for_for_asn_4753;
  wire CONVOLUTION_LOOP_for_for_for_asn_4755;
  wire CONVOLUTION_LOOP_for_for_for_asn_4757;
  wire CONVOLUTION_LOOP_for_for_for_asn_4759;
  wire CONVOLUTION_LOOP_for_for_for_asn_4761;
  wire CONVOLUTION_LOOP_for_for_for_asn_4763;
  wire CONVOLUTION_LOOP_for_for_for_asn_4765;
  wire CONVOLUTION_LOOP_for_for_for_asn_4767;
  wire CONVOLUTION_LOOP_for_for_for_asn_4769;
  wire CONVOLUTION_LOOP_for_for_for_asn_4771;
  wire CONVOLUTION_LOOP_for_for_for_asn_4773;
  wire CONVOLUTION_LOOP_for_for_for_asn_4775;
  wire CONVOLUTION_LOOP_for_for_for_asn_4777;
  wire CONVOLUTION_LOOP_for_for_for_asn_4779;
  wire CONVOLUTION_LOOP_for_for_for_asn_4781;
  wire CONVOLUTION_LOOP_for_for_for_asn_4783;
  wire CONVOLUTION_LOOP_for_for_for_asn_4785;
  wire CONVOLUTION_LOOP_for_for_for_asn_4787;
  wire CONVOLUTION_LOOP_for_for_for_asn_4789;
  wire CONVOLUTION_LOOP_for_for_for_asn_4791;
  wire CONVOLUTION_LOOP_for_for_for_asn_4793;
  wire CONVOLUTION_LOOP_for_for_for_asn_4795;
  wire CONVOLUTION_LOOP_for_for_for_asn_4797;
  wire CONVOLUTION_LOOP_for_for_for_asn_4799;
  wire CONVOLUTION_LOOP_for_for_for_asn_4801;
  wire CONVOLUTION_LOOP_for_for_for_asn_4803;
  wire CONVOLUTION_LOOP_for_for_for_asn_4805;
  wire CONVOLUTION_LOOP_for_for_for_asn_4807;
  wire CONVOLUTION_LOOP_for_for_for_asn_4809;
  wire CONVOLUTION_LOOP_for_for_for_asn_4811;
  wire CONVOLUTION_LOOP_for_for_for_asn_4813;
  wire CONVOLUTION_LOOP_for_for_for_asn_4815;
  wire CONVOLUTION_LOOP_for_for_for_asn_4817;
  wire CONVOLUTION_LOOP_for_for_for_asn_4819;
  wire CONVOLUTION_LOOP_for_for_for_asn_4821;
  wire CONVOLUTION_LOOP_for_for_for_asn_4823;
  wire CONVOLUTION_LOOP_for_for_for_asn_4825;
  wire CONVOLUTION_LOOP_for_for_for_asn_4827;
  wire CONVOLUTION_LOOP_for_for_for_asn_4829;
  wire CONVOLUTION_LOOP_for_for_for_asn_4831;
  wire CONVOLUTION_LOOP_for_for_for_asn_4833;
  wire CONVOLUTION_LOOP_for_for_for_asn_4835;
  wire CONVOLUTION_LOOP_for_for_for_asn_4837;
  wire CONVOLUTION_LOOP_for_for_for_asn_4839;
  wire CONVOLUTION_LOOP_for_for_for_asn_4841;
  wire CONVOLUTION_LOOP_for_for_for_asn_4843;
  wire CONVOLUTION_LOOP_for_for_for_asn_4845;
  wire CONVOLUTION_LOOP_for_for_for_asn_4847;
  wire CONVOLUTION_LOOP_for_for_for_asn_4849;
  wire CONVOLUTION_LOOP_for_for_for_asn_4851;
  wire CONVOLUTION_LOOP_for_for_for_asn_4853;
  wire CONVOLUTION_LOOP_for_for_for_asn_4855;
  wire CONVOLUTION_LOOP_for_for_for_asn_4857;
  wire CONVOLUTION_LOOP_for_for_for_asn_4859;
  wire CONVOLUTION_LOOP_for_for_for_asn_4861;
  wire CONVOLUTION_LOOP_for_for_for_asn_4863;
  wire CONVOLUTION_LOOP_for_for_for_asn_4865;
  wire CONVOLUTION_LOOP_for_for_for_asn_4867;
  wire CONVOLUTION_LOOP_for_for_for_asn_4869;
  wire CONVOLUTION_LOOP_for_for_for_asn_4871;
  wire CONVOLUTION_LOOP_for_for_for_asn_4873;
  wire CONVOLUTION_LOOP_for_for_for_asn_4875;
  wire CONVOLUTION_LOOP_for_for_for_asn_4877;
  wire CONVOLUTION_LOOP_for_for_for_asn_4879;
  wire CONVOLUTION_LOOP_for_for_for_asn_4881;
  wire CONVOLUTION_LOOP_for_for_for_asn_4883;
  wire CONVOLUTION_LOOP_for_for_for_asn_4885;
  wire CONVOLUTION_LOOP_for_for_for_asn_4887;
  wire CONVOLUTION_LOOP_for_for_for_asn_4889;
  wire CONVOLUTION_LOOP_for_for_for_asn_4891;
  wire CONVOLUTION_LOOP_for_for_for_asn_4893;
  wire CONVOLUTION_LOOP_for_for_for_asn_4895;
  wire CONVOLUTION_LOOP_for_for_for_asn_4897;
  wire CONVOLUTION_LOOP_for_for_for_asn_4899;
  wire CONVOLUTION_LOOP_for_for_for_asn_4901;
  wire CONVOLUTION_LOOP_for_for_for_asn_4903;
  wire CONVOLUTION_LOOP_for_for_for_asn_4905;
  wire CONVOLUTION_LOOP_for_for_for_asn_4907;
  wire CONVOLUTION_LOOP_for_for_for_asn_4909;
  wire CONVOLUTION_LOOP_for_for_for_asn_4911;
  wire CONVOLUTION_LOOP_for_for_for_asn_4913;
  wire CONVOLUTION_LOOP_for_for_for_asn_4915;
  wire CONVOLUTION_LOOP_for_for_for_asn_4917;
  wire CONVOLUTION_LOOP_for_for_for_asn_4919;
  wire CONVOLUTION_LOOP_for_for_for_asn_4921;
  wire CONVOLUTION_LOOP_for_for_for_asn_4923;
  wire CONVOLUTION_LOOP_for_for_for_asn_4925;
  wire CONVOLUTION_LOOP_for_for_for_asn_4927;
  wire CONVOLUTION_LOOP_for_for_for_asn_4929;
  wire CONVOLUTION_LOOP_for_for_for_asn_4931;
  wire CONVOLUTION_LOOP_for_for_for_asn_4933;
  wire CONVOLUTION_LOOP_for_for_for_asn_4935;
  wire CONVOLUTION_LOOP_for_for_for_asn_4937;
  wire CONVOLUTION_LOOP_for_for_for_asn_4939;
  wire CONVOLUTION_LOOP_for_for_for_asn_4941;
  wire CONVOLUTION_LOOP_for_for_for_asn_4943;
  wire CONVOLUTION_LOOP_for_for_for_asn_4945;
  wire CONVOLUTION_LOOP_for_for_for_asn_4947;
  wire CONVOLUTION_LOOP_for_for_for_asn_4949;
  wire CONVOLUTION_LOOP_for_for_for_asn_4951;
  wire CONVOLUTION_LOOP_for_for_for_asn_4953;
  wire CONVOLUTION_LOOP_for_for_for_asn_4955;
  wire CONVOLUTION_LOOP_for_for_for_asn_4957;
  wire CONVOLUTION_LOOP_for_for_for_asn_4959;
  wire CONVOLUTION_LOOP_for_for_for_asn_4961;
  wire CONVOLUTION_LOOP_for_for_for_asn_4963;
  wire CONVOLUTION_LOOP_for_for_for_asn_4965;
  wire CONVOLUTION_LOOP_for_for_for_asn_4967;
  wire CONVOLUTION_LOOP_for_for_for_asn_4969;
  wire CONVOLUTION_LOOP_for_for_for_asn_4971;
  wire CONVOLUTION_LOOP_for_for_for_asn_4973;
  wire CONVOLUTION_LOOP_for_for_for_asn_4975;
  wire CONVOLUTION_LOOP_for_for_for_asn_4977;
  wire CONVOLUTION_LOOP_for_for_for_asn_4979;
  wire CONVOLUTION_LOOP_for_for_for_asn_4981;
  wire CONVOLUTION_LOOP_for_for_for_asn_4983;
  wire CONVOLUTION_LOOP_for_for_for_asn_4985;
  wire CONVOLUTION_LOOP_for_for_for_asn_4987;
  wire CONVOLUTION_LOOP_for_for_for_asn_4989;
  wire CONVOLUTION_LOOP_for_for_for_asn_4991;
  wire CONVOLUTION_LOOP_for_for_for_asn_4993;
  wire CONVOLUTION_LOOP_for_for_for_asn_4995;
  wire CONVOLUTION_LOOP_for_for_for_asn_4997;
  wire CONVOLUTION_LOOP_for_for_for_asn_4999;
  wire CONVOLUTION_LOOP_for_for_for_asn_5001;
  wire CONVOLUTION_LOOP_for_for_for_asn_5003;
  wire CONVOLUTION_LOOP_for_for_for_asn_5005;
  wire CONVOLUTION_LOOP_for_for_for_asn_5007;
  wire CONVOLUTION_LOOP_for_for_for_asn_5009;
  wire CONVOLUTION_LOOP_for_for_for_asn_5011;
  wire CONVOLUTION_LOOP_for_for_for_asn_5013;
  wire CONVOLUTION_LOOP_for_for_for_asn_5015;
  wire CONVOLUTION_LOOP_for_for_for_asn_5017;
  wire CONVOLUTION_LOOP_for_for_for_asn_5019;
  wire CONVOLUTION_LOOP_for_for_for_asn_5021;
  wire CONVOLUTION_LOOP_for_for_for_asn_5023;
  wire CONVOLUTION_LOOP_for_for_for_asn_5025;
  wire CONVOLUTION_LOOP_for_for_for_asn_5027;
  wire CONVOLUTION_LOOP_for_for_for_asn_5029;
  wire CONVOLUTION_LOOP_for_for_for_asn_5031;
  wire CONVOLUTION_LOOP_for_for_for_asn_5033;
  wire CONVOLUTION_LOOP_for_for_for_asn_5035;
  wire CONVOLUTION_LOOP_for_for_for_asn_5037;
  wire CONVOLUTION_LOOP_for_for_for_asn_5039;
  wire CONVOLUTION_LOOP_for_for_for_asn_5041;
  wire CONVOLUTION_LOOP_for_for_for_asn_5043;
  wire CONVOLUTION_LOOP_for_for_for_asn_5045;
  wire CONVOLUTION_LOOP_for_for_for_asn_5047;
  wire CONVOLUTION_LOOP_for_for_for_asn_5049;
  wire CONVOLUTION_LOOP_for_for_for_asn_5051;
  wire CONVOLUTION_LOOP_for_for_for_asn_5053;
  wire CONVOLUTION_LOOP_for_for_for_asn_5055;
  wire CONVOLUTION_LOOP_for_for_for_asn_5057;
  wire CONVOLUTION_LOOP_for_for_for_asn_5059;
  wire CONVOLUTION_LOOP_for_for_for_asn_5061;
  wire CONVOLUTION_LOOP_for_for_for_asn_5063;
  wire CONVOLUTION_LOOP_for_for_for_asn_5065;
  wire CONVOLUTION_LOOP_for_for_for_asn_5067;
  wire CONVOLUTION_LOOP_for_for_for_asn_5069;
  wire CONVOLUTION_LOOP_for_for_for_asn_5071;
  wire CONVOLUTION_LOOP_for_for_for_asn_5073;
  wire CONVOLUTION_LOOP_for_for_for_asn_5075;
  wire CONVOLUTION_LOOP_for_for_for_asn_5077;
  wire CONVOLUTION_LOOP_for_for_for_asn_5079;
  wire CONVOLUTION_LOOP_for_for_for_asn_5081;
  wire CONVOLUTION_LOOP_for_for_for_asn_5083;
  wire CONVOLUTION_LOOP_for_for_for_asn_5085;
  wire CONVOLUTION_LOOP_for_for_for_asn_5087;
  wire CONVOLUTION_LOOP_for_for_for_asn_5089;
  wire CONVOLUTION_LOOP_for_for_for_asn_5091;
  wire CONVOLUTION_LOOP_for_for_for_asn_5093;
  wire CONVOLUTION_LOOP_for_for_for_asn_5095;
  wire CONVOLUTION_LOOP_for_for_for_asn_5097;
  wire CONVOLUTION_LOOP_for_for_for_asn_5099;
  wire CONVOLUTION_LOOP_for_for_for_asn_5101;
  wire CONVOLUTION_LOOP_for_for_for_asn_5103;
  wire CONVOLUTION_LOOP_for_for_for_asn_5105;
  wire CONVOLUTION_LOOP_for_for_for_asn_5107;
  wire CONVOLUTION_LOOP_for_for_for_asn_5109;
  wire CONVOLUTION_LOOP_for_for_for_asn_5111;
  wire CONVOLUTION_LOOP_for_for_for_asn_5113;
  wire CONVOLUTION_LOOP_for_for_for_asn_5115;
  wire CONVOLUTION_LOOP_for_for_for_asn_5117;
  wire CONVOLUTION_LOOP_for_for_for_asn_5119;
  wire CONVOLUTION_LOOP_for_for_for_asn_5121;
  wire CONVOLUTION_LOOP_for_for_for_asn_5123;
  wire CONVOLUTION_LOOP_for_for_for_asn_5125;
  wire CONVOLUTION_LOOP_for_for_for_asn_5127;
  wire CONVOLUTION_LOOP_for_for_for_asn_5129;
  wire CONVOLUTION_LOOP_for_for_for_asn_5131;
  wire CONVOLUTION_LOOP_for_for_for_asn_5133;
  wire CONVOLUTION_LOOP_for_for_for_asn_5135;
  wire CONVOLUTION_LOOP_for_for_for_asn_5137;
  wire CONVOLUTION_LOOP_for_for_for_asn_5139;
  wire CONVOLUTION_LOOP_for_for_for_asn_5141;
  wire CONVOLUTION_LOOP_for_for_for_asn_5143;
  wire CONVOLUTION_LOOP_for_for_for_asn_5145;
  wire CONVOLUTION_LOOP_for_for_for_asn_5147;
  wire CONVOLUTION_LOOP_for_for_for_asn_5149;
  wire CONVOLUTION_LOOP_for_for_for_asn_5151;
  wire CONVOLUTION_LOOP_for_for_for_asn_5153;
  wire CONVOLUTION_LOOP_for_for_for_asn_5155;
  wire CONVOLUTION_LOOP_for_for_for_asn_5157;
  wire CONVOLUTION_LOOP_for_for_for_asn_5159;
  wire CONVOLUTION_LOOP_for_for_for_asn_5161;
  wire CONVOLUTION_LOOP_for_for_for_asn_5163;
  wire CONVOLUTION_LOOP_for_for_for_asn_5165;
  wire CONVOLUTION_LOOP_for_for_for_asn_5167;
  wire CONVOLUTION_LOOP_for_for_for_asn_5169;
  wire CONVOLUTION_LOOP_for_for_for_asn_5171;
  wire CONVOLUTION_LOOP_for_for_for_asn_5173;
  wire CONVOLUTION_LOOP_for_for_for_asn_5175;
  wire CONVOLUTION_LOOP_for_for_for_asn_5177;
  wire CONVOLUTION_LOOP_for_for_for_asn_5179;
  wire CONVOLUTION_LOOP_for_for_for_asn_5181;
  wire CONVOLUTION_LOOP_for_for_for_asn_5183;
  wire CONVOLUTION_LOOP_for_for_for_asn_5185;
  wire CONVOLUTION_LOOP_for_for_for_asn_5187;
  wire CONVOLUTION_LOOP_for_for_for_asn_5189;
  wire CONVOLUTION_LOOP_for_for_for_asn_5191;
  wire CONVOLUTION_LOOP_for_for_for_asn_5193;
  wire CONVOLUTION_LOOP_for_for_for_asn_5195;
  wire CONVOLUTION_LOOP_for_for_for_asn_5197;
  wire CONVOLUTION_LOOP_for_for_for_asn_5199;
  wire CONVOLUTION_LOOP_for_for_for_asn_5201;
  wire CONVOLUTION_LOOP_for_for_for_asn_5203;
  wire CONVOLUTION_LOOP_for_for_for_asn_5205;
  wire CONVOLUTION_LOOP_for_for_for_asn_5207;
  wire CONVOLUTION_LOOP_for_for_for_asn_5209;
  wire CONVOLUTION_LOOP_for_for_for_asn_5211;
  wire CONVOLUTION_LOOP_for_for_for_asn_5213;
  wire CONVOLUTION_LOOP_for_for_for_asn_5215;
  wire CONVOLUTION_LOOP_for_for_for_asn_5217;
  wire CONVOLUTION_LOOP_for_for_for_asn_5219;
  wire CONVOLUTION_LOOP_for_for_for_asn_5221;
  wire CONVOLUTION_LOOP_for_for_for_asn_5223;
  wire CONVOLUTION_LOOP_for_for_for_asn_5225;
  wire CONVOLUTION_LOOP_for_for_for_asn_5227;
  wire CONVOLUTION_LOOP_for_for_for_asn_5229;
  wire CONVOLUTION_LOOP_for_for_for_asn_5231;
  wire CONVOLUTION_LOOP_for_for_for_asn_5233;
  wire CONVOLUTION_LOOP_for_for_for_asn_5235;
  wire CONVOLUTION_LOOP_for_for_for_asn_5237;
  wire CONVOLUTION_LOOP_for_for_for_asn_5239;
  wire CONVOLUTION_LOOP_for_for_for_asn_5241;
  wire CONVOLUTION_LOOP_for_for_for_asn_5243;
  wire CONVOLUTION_LOOP_for_for_for_asn_5245;
  wire CONVOLUTION_LOOP_for_for_for_asn_5247;
  wire CONVOLUTION_LOOP_for_for_for_asn_5249;
  wire CONVOLUTION_LOOP_for_for_for_asn_5251;
  wire CONVOLUTION_LOOP_for_for_for_asn_5253;
  wire CONVOLUTION_LOOP_for_for_for_asn_5255;
  wire CONVOLUTION_LOOP_for_for_for_asn_5257;
  wire CONVOLUTION_LOOP_for_for_for_asn_5259;
  wire CONVOLUTION_LOOP_for_for_for_asn_5261;
  wire CONVOLUTION_LOOP_for_for_for_asn_5263;
  wire CONVOLUTION_LOOP_for_for_for_asn_5265;
  wire CONVOLUTION_LOOP_for_for_for_asn_5267;
  wire CONVOLUTION_LOOP_for_for_for_asn_5269;
  wire CONVOLUTION_LOOP_for_for_for_asn_5271;
  wire CONVOLUTION_LOOP_for_for_for_asn_5273;
  wire CONVOLUTION_LOOP_for_for_for_asn_5275;
  wire CONVOLUTION_LOOP_for_for_for_asn_5277;
  wire CONVOLUTION_LOOP_for_for_for_asn_5279;
  wire CONVOLUTION_LOOP_for_for_for_asn_5281;
  wire CONVOLUTION_LOOP_for_for_for_asn_5283;
  wire CONVOLUTION_LOOP_for_for_for_asn_5285;
  wire CONVOLUTION_LOOP_for_for_for_asn_5287;
  wire CONVOLUTION_LOOP_for_for_for_asn_5289;
  wire CONVOLUTION_LOOP_for_for_for_asn_5291;
  wire CONVOLUTION_LOOP_for_for_for_asn_5293;
  wire CONVOLUTION_LOOP_for_for_for_asn_5295;
  wire CONVOLUTION_LOOP_for_for_for_asn_5297;
  wire CONVOLUTION_LOOP_for_for_for_asn_5299;
  wire CONVOLUTION_LOOP_for_for_for_asn_5301;
  wire CONVOLUTION_LOOP_for_for_for_asn_5303;
  wire CONVOLUTION_LOOP_for_for_for_asn_5305;
  wire CONVOLUTION_LOOP_for_for_for_asn_5307;
  wire CONVOLUTION_LOOP_for_for_for_asn_5309;
  wire CONVOLUTION_LOOP_for_for_for_asn_5311;
  wire CONVOLUTION_LOOP_for_for_for_asn_5313;
  wire CONVOLUTION_LOOP_for_for_for_asn_5315;
  wire CONVOLUTION_LOOP_for_for_for_asn_5317;
  wire CONVOLUTION_LOOP_for_for_for_asn_5319;
  wire CONVOLUTION_LOOP_for_for_for_asn_5321;
  wire CONVOLUTION_LOOP_for_for_for_asn_5323;
  wire CONVOLUTION_LOOP_for_for_for_asn_5325;
  wire CONVOLUTION_LOOP_for_for_for_asn_5327;
  wire CONVOLUTION_LOOP_for_for_for_asn_5329;
  wire CONVOLUTION_LOOP_for_for_for_asn_5331;
  wire CONVOLUTION_LOOP_for_for_for_asn_5333;
  wire CONVOLUTION_LOOP_for_for_for_asn_5335;
  wire CONVOLUTION_LOOP_for_for_for_asn_5337;
  wire CONVOLUTION_LOOP_for_for_for_asn_5339;
  wire CONVOLUTION_LOOP_for_for_for_asn_5341;
  wire CONVOLUTION_LOOP_for_for_for_asn_5343;
  wire CONVOLUTION_LOOP_for_for_for_asn_5345;
  wire CONVOLUTION_LOOP_for_for_for_asn_5347;
  wire CONVOLUTION_LOOP_for_for_for_asn_5349;
  wire CONVOLUTION_LOOP_for_for_for_asn_5351;
  wire CONVOLUTION_LOOP_for_for_for_asn_5353;
  wire CONVOLUTION_LOOP_for_for_for_asn_5355;
  wire CONVOLUTION_LOOP_for_for_for_asn_5357;
  wire CONVOLUTION_LOOP_for_for_for_asn_5359;
  wire CONVOLUTION_LOOP_for_for_for_asn_5361;
  wire CONVOLUTION_LOOP_for_for_for_asn_5363;
  wire CONVOLUTION_LOOP_for_for_for_asn_5365;
  wire CONVOLUTION_LOOP_for_for_for_asn_5367;
  wire CONVOLUTION_LOOP_for_for_for_asn_5369;
  wire CONVOLUTION_LOOP_for_for_for_asn_5371;
  wire CONVOLUTION_LOOP_for_for_for_asn_5373;
  wire CONVOLUTION_LOOP_for_for_for_asn_5375;
  wire CONVOLUTION_LOOP_for_for_for_asn_5377;
  wire CONVOLUTION_LOOP_for_for_for_asn_5379;
  wire CONVOLUTION_LOOP_for_for_for_asn_5381;
  wire CONVOLUTION_LOOP_for_for_for_asn_5383;
  wire CONVOLUTION_LOOP_for_for_for_asn_5385;
  wire CONVOLUTION_LOOP_for_for_for_asn_5387;
  wire CONVOLUTION_LOOP_for_for_for_asn_5389;
  wire CONVOLUTION_LOOP_for_for_for_asn_5391;
  wire CONVOLUTION_LOOP_for_for_for_asn_5393;
  wire CONVOLUTION_LOOP_for_for_for_asn_5395;
  wire CONVOLUTION_LOOP_for_for_for_asn_5397;
  wire CONVOLUTION_LOOP_for_for_for_asn_5399;
  wire CONVOLUTION_LOOP_for_for_for_asn_5401;
  wire CONVOLUTION_LOOP_for_for_for_asn_5403;
  wire CONVOLUTION_LOOP_for_for_for_asn_5405;
  wire CONVOLUTION_LOOP_for_for_for_asn_5407;
  wire CONVOLUTION_LOOP_for_for_for_asn_5409;
  wire CONVOLUTION_LOOP_for_for_for_asn_5411;
  wire CONVOLUTION_LOOP_for_for_for_asn_5413;
  wire CONVOLUTION_LOOP_for_for_for_asn_5415;
  wire CONVOLUTION_LOOP_for_for_for_asn_5417;
  wire CONVOLUTION_LOOP_for_for_for_asn_5419;
  wire CONVOLUTION_LOOP_for_for_for_asn_5421;
  wire CONVOLUTION_LOOP_for_for_for_asn_5423;
  wire CONVOLUTION_LOOP_for_for_for_asn_5425;
  wire CONVOLUTION_LOOP_for_for_for_asn_5427;
  wire CONVOLUTION_LOOP_for_for_for_asn_5429;
  wire CONVOLUTION_LOOP_for_for_for_asn_5431;
  wire CONVOLUTION_LOOP_for_for_for_asn_5433;
  wire CONVOLUTION_LOOP_for_for_for_asn_5435;
  wire CONVOLUTION_LOOP_for_for_for_asn_5437;
  wire CONVOLUTION_LOOP_for_for_for_asn_5439;
  wire CONVOLUTION_LOOP_for_for_for_asn_5441;
  wire CONVOLUTION_LOOP_for_for_for_asn_5443;
  wire CONVOLUTION_LOOP_for_for_for_asn_5445;
  wire CONVOLUTION_LOOP_for_for_for_asn_5447;
  wire CONVOLUTION_LOOP_for_for_for_asn_5449;
  wire CONVOLUTION_LOOP_for_for_for_asn_5451;
  wire CONVOLUTION_LOOP_for_for_for_asn_5453;
  wire CONVOLUTION_LOOP_for_for_for_asn_5455;
  wire CONVOLUTION_LOOP_for_for_for_asn_5457;
  wire CONVOLUTION_LOOP_for_for_for_asn_5459;
  wire CONVOLUTION_LOOP_for_for_for_asn_5461;
  wire CONVOLUTION_LOOP_for_for_for_asn_5463;
  wire CONVOLUTION_LOOP_for_for_for_asn_5465;
  wire CONVOLUTION_LOOP_for_for_for_asn_5467;
  wire CONVOLUTION_LOOP_for_for_for_asn_5469;
  wire CONVOLUTION_LOOP_for_for_for_asn_5471;
  wire CONVOLUTION_LOOP_for_for_for_asn_5473;
  wire CONVOLUTION_LOOP_for_for_for_asn_5475;
  wire CONVOLUTION_LOOP_for_for_for_asn_5477;
  wire CONVOLUTION_LOOP_for_for_for_asn_5479;
  wire CONVOLUTION_LOOP_for_for_for_asn_5481;
  wire CONVOLUTION_LOOP_for_for_for_asn_5483;
  wire CONVOLUTION_LOOP_for_for_for_asn_5485;
  wire CONVOLUTION_LOOP_for_for_for_asn_5487;
  wire CONVOLUTION_LOOP_for_for_for_asn_5489;
  wire CONVOLUTION_LOOP_for_for_for_asn_5491;
  wire CONVOLUTION_LOOP_for_for_for_asn_5493;
  wire CONVOLUTION_LOOP_for_for_for_asn_5495;
  wire CONVOLUTION_LOOP_for_for_for_asn_5497;
  wire CONVOLUTION_LOOP_for_for_for_asn_5499;
  wire CONVOLUTION_LOOP_for_for_for_asn_5501;
  wire CONVOLUTION_LOOP_for_for_for_asn_5503;
  wire CONVOLUTION_LOOP_for_for_for_asn_5505;
  wire CONVOLUTION_LOOP_for_for_for_asn_5507;
  wire CONVOLUTION_LOOP_for_for_for_asn_5509;
  wire CONVOLUTION_LOOP_for_for_for_asn_5511;
  wire CONVOLUTION_LOOP_for_for_for_asn_5513;
  wire CONVOLUTION_LOOP_for_for_for_asn_5515;
  wire CONVOLUTION_LOOP_for_for_for_asn_5517;
  wire COMPUTE_LOOP_asn_44;
  wire COMPUTE_LOOP_asn_46;
  wire CONVOLUTION_LOOP_for_and_3_rgt;
  wire CONVOLUTION_LOOP_for_and_4_rgt;
  wire and_88_rgt;
  wire CONVOLUTION_LOOP_for_for_and_3_rgt;
  wire CONVOLUTION_LOOP_for_for_and_4_rgt;
  wire and_90_rgt;
  wire CONVOLUTION_LOOP_for_for_for_and_2588_rgt;
  wire CONVOLUTION_LOOP_for_for_for_and_2589_rgt;
  wire CONVOLUTION_LOOP_for_for_for_y_and_rgt;
  wire CONVOLUTION_LOOP_for_for_for_y_and_1_rgt;
  wire CONVOLUTION_LOOP_for_for_for_j_and_cse;
  reg [4:0] reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse;
  reg [2:0] reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse;
  wire CONVOLUTION_LOOP_for_for_for_for_for_n_and_itm;
  wire CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm;
  wire operator_8_false_3_acc_itm_4_1;
  wire operator_8_false_4_acc_itm_4;
  wire operator_8_false_5_acc_itm_3_1;
  wire operator_8_false_6_acc_itm_3_1;

  wire[0:0] mux_37_nl;
  wire[0:0] or_89_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl;
  wire[29:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_nl;
  wire[29:0] CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_2_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_12_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_24_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_36_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_48_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_60_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_72_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_84_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_96_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_108_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_120_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_132_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_144_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_156_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_168_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_180_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_192_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_204_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_216_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_228_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_240_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_252_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_264_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_276_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_288_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_300_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_312_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_324_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_336_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_348_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_360_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_372_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_384_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_396_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_408_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_420_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_432_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_444_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_456_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_468_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_480_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_492_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_504_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_516_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_528_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_540_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_552_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_564_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_576_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_588_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_600_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_612_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_624_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_636_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_648_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_660_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_672_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_684_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_696_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_708_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_720_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_732_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_744_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_756_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_768_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_780_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_792_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_804_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_816_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_828_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_840_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_852_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_864_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_876_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_888_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_900_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_912_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_924_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_936_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_948_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_960_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_972_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_984_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_996_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1008_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1020_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1032_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1044_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1056_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1068_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1080_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1092_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1104_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1116_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1128_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1140_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1152_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1164_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1176_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1188_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1200_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1212_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1224_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1236_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1248_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1260_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1272_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1284_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1296_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1308_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1320_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1332_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1344_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1356_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1368_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1380_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1392_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1404_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1416_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1428_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1440_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1452_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1464_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1476_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1488_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1500_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1512_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1524_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1536_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1548_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1560_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1572_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1584_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1596_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1608_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1620_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1632_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1644_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1656_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1668_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1680_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1692_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1704_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1716_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1728_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1740_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1752_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1764_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1776_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1788_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1800_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1812_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1824_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1836_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1848_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1860_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1872_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1884_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1896_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1908_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1920_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1932_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1944_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1938_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1926_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1914_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1902_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1890_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1878_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1866_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1854_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1842_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1830_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1818_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1806_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1794_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1782_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1770_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1758_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1746_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1734_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1722_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1710_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1698_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1686_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1674_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1662_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1650_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1638_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1626_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1614_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1602_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1590_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1578_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1566_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1554_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1542_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1530_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1518_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1506_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1494_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1482_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1470_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1458_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1446_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1434_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1422_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1410_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1398_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1386_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1374_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1362_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1350_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1338_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1326_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1314_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1302_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1290_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1278_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1266_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1254_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1242_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1230_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1218_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1206_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1194_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1182_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1170_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1158_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1146_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1134_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1122_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1110_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1098_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1086_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1074_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1062_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1050_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1038_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1026_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1014_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_1002_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_990_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_978_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_966_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_954_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_942_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_930_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_918_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_906_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_894_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_882_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_870_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_858_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_846_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_834_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_822_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_810_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_798_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_786_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_774_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_762_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_750_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_738_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_726_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_714_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_702_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_690_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_678_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_666_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_654_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_642_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_630_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_618_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_606_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_594_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_582_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_570_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_558_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_546_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_534_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_522_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_510_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_498_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_486_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_474_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_462_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_450_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_438_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_426_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_414_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_402_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_390_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_378_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_366_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_354_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_342_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_330_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_318_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_306_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_294_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_282_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_270_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_258_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_246_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_234_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_222_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_210_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_198_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_186_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_174_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_162_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_150_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_138_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_126_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_114_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_102_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_90_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_78_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_66_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_54_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_42_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_30_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_18_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_mux_6_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_10_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_22_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_34_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_46_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_58_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_70_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_82_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_94_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_106_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_118_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_130_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_142_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_154_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_166_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_178_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_190_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_202_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_214_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_226_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_238_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_250_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_262_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_274_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_286_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_298_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_310_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_322_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_334_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_346_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_358_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_370_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_382_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_394_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_406_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_418_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_430_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_442_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_454_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_466_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_478_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_490_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_502_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_514_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_526_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_538_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_550_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_562_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_574_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_586_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_598_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_610_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_622_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_634_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_646_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_658_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_670_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_682_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_694_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_706_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_718_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_730_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_742_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_754_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_766_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_778_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_790_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_802_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_814_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_826_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_838_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_850_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_862_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_874_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_886_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_898_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_910_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_922_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_934_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_946_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_958_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_970_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_982_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_994_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1006_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1018_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1030_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1042_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1054_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1066_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1078_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1090_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1102_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1114_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1126_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1138_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1150_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1162_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1174_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1186_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1198_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1210_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1222_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1234_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1246_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1258_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1270_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1282_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1294_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1306_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1318_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1330_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1342_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1354_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1366_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1378_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1390_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1402_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1414_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1426_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1438_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1450_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1462_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1474_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1486_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1498_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1510_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1522_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1534_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1546_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1558_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1570_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1582_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1594_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1606_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1618_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1630_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1642_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1654_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1666_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1678_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1690_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1702_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1714_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1726_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1738_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1750_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1762_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1774_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1786_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1798_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1810_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1822_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1834_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1846_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1858_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1870_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1882_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1894_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1906_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1918_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1930_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1942_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1936_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1924_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1912_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1900_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1888_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1876_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1864_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1852_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1840_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1828_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1816_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1804_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1792_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1780_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1768_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1756_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1744_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1732_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1720_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1708_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1696_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1684_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1672_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1660_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1648_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1636_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1624_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1612_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1600_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1588_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1576_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1564_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1552_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1540_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1528_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1516_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1504_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1492_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1480_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1468_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1456_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1444_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1432_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1420_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1408_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1396_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1384_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1372_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1360_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1348_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1336_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1324_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1312_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1300_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1288_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1276_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1264_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1252_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1240_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1228_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1216_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1204_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1192_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1180_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1168_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1156_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1144_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1132_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1120_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1108_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1096_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1084_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1072_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1060_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1048_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1036_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1024_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1012_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_1000_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_988_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_976_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_964_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_952_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_940_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_928_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_916_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_904_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_892_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_880_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_868_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_856_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_844_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_832_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_820_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_808_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_796_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_784_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_772_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_760_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_748_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_736_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_724_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_712_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_700_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_688_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_676_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_664_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_652_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_640_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_628_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_616_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_604_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_592_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_580_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_568_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_556_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_544_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_532_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_520_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_508_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_496_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_484_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_472_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_460_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_448_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_436_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_424_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_412_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_400_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_388_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_376_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_364_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_352_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_340_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_328_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_316_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_304_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_292_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_280_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_268_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_256_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_244_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_232_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_220_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_208_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_196_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_184_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_172_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_160_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_148_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_136_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_124_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_112_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_100_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_88_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_76_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_64_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_52_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_40_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_28_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_16_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_mux_4_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_8_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_20_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_32_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_44_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_56_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_68_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_80_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_92_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_308_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_320_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_332_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_344_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_356_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_368_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_380_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_392_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_404_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_416_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_428_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_440_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_452_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_464_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_476_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_488_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_500_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_512_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_524_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_536_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_548_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_560_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_572_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_584_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_596_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_608_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_620_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_632_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_644_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_656_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_668_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_680_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_692_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_704_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_716_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_728_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_740_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_752_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_764_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_776_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_788_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_800_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_812_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_824_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_836_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_848_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_860_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_872_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_884_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_896_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_908_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_920_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_932_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_944_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_956_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_968_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1304_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1316_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1328_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1340_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1352_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1364_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1376_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1388_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1400_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1412_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1424_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1436_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1448_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1460_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1472_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1484_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1496_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1508_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1520_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1532_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1544_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1556_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1568_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1580_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1592_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1604_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1616_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1628_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1640_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1652_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1664_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1676_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1688_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1700_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1712_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1724_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1736_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1748_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1760_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1772_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1784_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1796_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1808_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1820_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1832_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1844_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1856_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1868_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1880_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1892_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1904_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1916_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1928_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1940_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1934_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1922_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1910_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1898_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1886_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1874_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1862_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1850_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1838_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1826_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1814_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1802_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1790_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1778_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1766_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1754_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1742_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1730_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1718_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1706_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1694_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1682_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1670_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1658_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1646_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1634_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1622_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1610_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1598_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1586_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1574_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1562_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1550_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1538_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1526_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1514_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1502_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1478_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1466_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1454_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1442_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1430_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1418_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1406_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1394_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1382_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1370_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1358_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1346_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1334_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_962_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_950_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_938_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_926_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_914_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_902_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_890_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_878_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_866_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_854_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_842_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_830_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_818_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_806_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_794_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_782_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_770_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_758_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_746_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_734_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_722_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_710_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_698_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_686_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_674_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_662_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_650_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_638_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_626_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_614_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_602_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_590_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_578_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_566_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_554_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_542_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_530_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_518_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_506_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_494_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_482_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_470_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_458_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_446_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_434_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_422_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_410_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_398_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_386_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_374_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_362_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_350_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_338_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_326_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_98_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_86_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_74_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_62_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_50_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_38_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_26_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_14_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_2_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_acc_mux_5_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_acc_mux_3_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_not_28_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_acc_mux_1_nl;
  wire[2:0] CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_and_nl;
  wire[0:0] or_277_nl;
  wire[0:0] and_74_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] nor_51_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl;
  wire[14:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl;
  wire[15:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl;
  wire[18:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl;
  wire[15:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl;
  wire[16:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl;
  wire[20:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl;
  wire[12:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_4_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl;
  wire[11:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl;
  wire[10:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_5_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_nl;
  wire[23:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_nl;
  wire[15:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_1_nl;
  wire[20:0] nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_1_nl;
  wire[12:0] CONVOLUTION_LOOP_for_for_for_for_for_mul_2_nl;
  wire[0:0] and_84_nl;
  wire[12:0] CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl;
  wire[13:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl;
  wire[12:0] CONVOLUTION_LOOP_for_for_for_index_out_mul_2_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_index_out_mul_nl;
  wire[18:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_nl;
  wire[13:0] CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl;
  wire[15:0] nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl;
  wire[0:0] CONVOLUTION_LOOP_CONVOLUTION_LOOP_CONVOLUTION_LOOP_COMPUTE_LOOP_not_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_mux_1954_nl;
  wire[0:0] CONVOLUTION_LOOP_mux_6_nl;
  wire[7:0] if_acc_nl;
  wire[8:0] nl_if_acc_nl;
  wire[7:0] operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_acc_nl;
  wire[0:0] operator_42_true_and_nl;
  wire[7:0] if_acc_6_nl;
  wire[8:0] nl_if_acc_6_nl;
  wire[7:0] operator_43_true_1_acc_nl;
  wire[8:0] nl_operator_43_true_1_acc_nl;
  wire[0:0] operator_42_true_1_and_nl;
  wire[0:0] COMPUTE_LOOP_mux_4_nl;
  wire[0:0] CONVOLUTION_LOOP_for_mux_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_mux_1_nl;
  wire[44:0] CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl;
  wire[6:0] n_w_in_acc_nl;
  wire[7:0] nl_n_w_in_acc_nl;
  wire[6:0] n_h_in_acc_nl;
  wire[7:0] nl_n_h_in_acc_nl;
  wire[54:0] CONVOLUTION_LOOP_for_for_for_else_nor_1_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_974_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_978_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_975_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_976_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_977_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_984_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_978_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_979_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_988_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_980_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_981_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_982_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_983_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_996_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_984_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_985_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_986_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_987_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_988_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_989_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_990_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_991_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_992_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_993_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_994_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_995_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_996_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_997_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_998_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_999_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_if_mux_1297_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_for_and_7_nl;
  wire[7:0] operator_43_true_operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_operator_43_true_acc_nl;
  wire[0:0] operator_43_true_and_nl;
  wire[8:0] pad_acc_2_nl;
  wire[9:0] nl_pad_acc_2_nl;
  wire[16:0] pad_mul_nl;
  wire signed [17:0] nl_pad_mul_nl;
  wire[8:0] operator_8_false_acc_nl;
  wire[9:0] nl_operator_8_false_acc_nl;
  wire[0:0] COMPUTE_LOOP_not_35_nl;
  wire[0:0] CONVOLUTION_LOOP_not_13_nl;
  wire[4:0] operator_8_false_3_acc_nl;
  wire[5:0] nl_operator_8_false_3_acc_nl;
  wire[4:0] operator_8_false_4_acc_nl;
  wire[5:0] nl_operator_8_false_4_acc_nl;
  wire[3:0] operator_8_false_5_acc_nl;
  wire[4:0] nl_operator_8_false_5_acc_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_not_24_nl;
  wire[0:0] CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_4_nl;
  wire[7:0] CONVOLUTION_LOOP_for_for_for_x_mul_nl;
  wire[12:0] nl_CONVOLUTION_LOOP_for_for_for_x_mul_nl;
  wire[0:0] and_17_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] or_81_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] or_87_nl;
  wire[3:0] operator_8_false_6_acc_nl;
  wire[4:0] nl_operator_8_false_6_acc_nl;
  wire[7:0] CONVOLUTION_LOOP_for_for_for_for_for_mux_6_nl;
  wire[0:0] and_275_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_compute_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg;
  assign nl_compute_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg = and_dcpl_7
      & (fsm_output[1]);
  wire [0:0] nl_compute_core_plm_outputs_rsci_1_inst_plm_outputs_rsci_oswt_unreg;
  assign nl_compute_core_plm_outputs_rsci_1_inst_plm_outputs_rsci_oswt_unreg = and_dcpl_28
      & plm_outputs_rsci_bawt & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_3 & main_stage_v_3;
  wire [0:0] nl_compute_core_plm_outputs_rsc_rls_obj_inst_plm_outputs_rsc_rls_obj_oswt_unreg;
  assign nl_compute_core_plm_outputs_rsc_rls_obj_inst_plm_outputs_rsc_rls_obj_oswt_unreg
      = or_dcpl_16 & or_dcpl_14 & plm_outputs_rsc_rls_obj_bawt & exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_3
      & main_stage_v_3;
  esp_acc_conv2d_cxx_catapult_compute_core_conf_info_rsci compute_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(nl_compute_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg[0:0]),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_iswt0(reg_conf_info_rsci_iswt0_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsci_1 compute_core_plm_inputs_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsci_q_d(plm_inputs_rsci_q_d),
      .plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsci_oswt_unreg(or_tmp_109),
      .plm_inputs_rsci_bawt(plm_inputs_rsci_bawt),
      .plm_inputs_rsci_iswt0(reg_plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .plm_inputs_rsci_q_d_mxwt(plm_inputs_rsci_q_d_mxwt),
      .plm_inputs_rsci_iswt0_pff(or_tmp_108)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsci_1 compute_core_plm_filters_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsci_q_d(plm_filters_rsci_q_d),
      .plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsci_oswt_unreg(or_tmp_109),
      .plm_filters_rsci_bawt(plm_filters_rsci_bawt),
      .plm_filters_rsci_iswt0(reg_plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .plm_filters_rsci_q_d_mxwt(plm_filters_rsci_q_d_mxwt),
      .plm_filters_rsci_iswt0_pff(or_tmp_108)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsci_1 compute_core_plm_outputs_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsci_oswt_unreg(nl_compute_core_plm_outputs_rsci_1_inst_plm_outputs_rsci_oswt_unreg[0:0]),
      .plm_outputs_rsci_bawt(plm_outputs_rsci_bawt),
      .plm_outputs_rsci_iswt0(reg_plm_outputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse),
      .plm_outputs_rsci_we_d_pff(plm_outputs_rsci_we_d_iff),
      .plm_outputs_rsci_iswt0_pff(and_50_rmff)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_done_rsci compute_core_done_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(and_dcpl_32),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_iswt0(reg_done_rsci_ivld_core_psct_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_rls_obj compute_core_plm_outputs_rsc_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_rls_lz(plm_outputs_rsc_rls_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsc_rls_obj_oswt_unreg(nl_compute_core_plm_outputs_rsc_rls_obj_inst_plm_outputs_rsc_rls_obj_oswt_unreg[0:0]),
      .plm_outputs_rsc_rls_obj_bawt(plm_outputs_rsc_rls_obj_bawt),
      .plm_outputs_rsc_rls_obj_iswt0(reg_plm_filters_rsc_rls_obj_oswt_cse)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_rls_obj compute_core_plm_inputs_rsc_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_rls_lz(plm_inputs_rsc_rls_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_inputs_rsc_rls_obj_oswt_unreg(and_34_rmff),
      .plm_inputs_rsc_rls_obj_bawt(plm_inputs_rsc_rls_obj_bawt),
      .plm_inputs_rsc_rls_obj_iswt0(reg_plm_filters_rsc_rls_obj_ld_core_psct_cse)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_rls_obj compute_core_plm_filters_rsc_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_rls_lz(plm_filters_rsc_rls_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_filters_rsc_rls_obj_oswt_unreg(and_34_rmff),
      .plm_filters_rsc_rls_obj_bawt(plm_filters_rsc_rls_obj_bawt),
      .plm_filters_rsc_rls_obj_iswt0(reg_plm_filters_rsc_rls_obj_ld_core_psct_cse)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_filters_rsc_req_obj compute_core_plm_filters_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_req_vz(plm_filters_rsc_req_vz),
      .core_wen(core_wen),
      .plm_filters_rsc_req_obj_oswt_unreg(and_235_cse),
      .plm_filters_rsc_req_obj_bawt(plm_filters_rsc_req_obj_bawt),
      .plm_filters_rsc_req_obj_iswt0(plm_filters_rsc_req_obj_iswt0),
      .plm_filters_rsc_req_obj_wen_comp(plm_filters_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_inputs_rsc_req_obj compute_core_plm_inputs_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_inputs_rsc_req_vz(plm_inputs_rsc_req_vz),
      .core_wen(core_wen),
      .plm_inputs_rsc_req_obj_oswt_unreg(and_235_cse),
      .plm_inputs_rsc_req_obj_bawt(plm_inputs_rsc_req_obj_bawt),
      .plm_inputs_rsc_req_obj_iswt0(plm_inputs_rsc_req_obj_iswt0),
      .plm_inputs_rsc_req_obj_wen_comp(plm_inputs_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_plm_outputs_rsc_req_obj compute_core_plm_outputs_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_req_vz(plm_outputs_rsc_req_vz),
      .core_wen(core_wen),
      .plm_outputs_rsc_req_obj_oswt_unreg(and_dcpl_11),
      .plm_outputs_rsc_req_obj_bawt(plm_outputs_rsc_req_obj_bawt),
      .plm_outputs_rsc_req_obj_iswt0(plm_outputs_rsc_req_obj_iswt0),
      .plm_outputs_rsc_req_obj_wen_comp(plm_outputs_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_staller compute_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .plm_filters_rsc_req_obj_wen_comp(plm_filters_rsc_req_obj_wen_comp),
      .plm_inputs_rsc_req_obj_wen_comp(plm_inputs_rsc_req_obj_wen_comp),
      .plm_outputs_rsc_req_obj_wen_comp(plm_outputs_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_compute_core_core_fsm compute_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign or_113_cse = (~((operator_8_false_7_acc_tmp[8]) | CONVOLUTION_LOOP_if_CONVOLUTION_LOOP_if_nand_tmp))
      | (CONVOLUTION_LOOP_acc_tmp[5]);
  assign COMPUTE_LOOP_and_cse = core_wen & (~((~ and_9_tmp) | (fsm_output[0])));
  assign and_235_cse = exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_1 & and_7_tmp;
  assign and_34_rmff = and_5_tmp & exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_2;
  assign and_50_rmff = exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_2 & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2
      & and_5_tmp;
  assign CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff = MUX_v_14_2_2(CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2,
      plm_outputs_rsci_wadr_d_reg, or_dcpl_22);
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl = MUX_s_1_324_2(COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_1_mx0, COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_1_mx0, {reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse
      , reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0});
  assign CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_1_nl
      = ~((~(CONVOLUTION_LOOP_for_for_for_if_1_mux_2_nl | CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1))
      | CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_rmff = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_1_nl,
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5,
      or_dcpl_22);
  assign CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl = ~(MUX_v_30_2_2((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_45_1_1[29:0]),
      30'b111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_nl
      = ~(MUX_v_30_2_2(CONVOLUTION_LOOP_for_for_for_if_1_nor_3_nl, 30'b111111111111111111111111111111,
      CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff = MUX_v_30_2_2(CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_nl,
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4,
      or_dcpl_22);
  assign CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_2_nl
      = ~((~((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_45_1_1[30])
      | CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_2_nl,
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3,
      or_dcpl_22);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff = MUX_v_16_2_2(CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1,
      plm_filters_rsci_radr_d_reg, or_tmp_111);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff = MUX_v_14_2_2(CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1,
      plm_inputs_rsci_radr_d_reg, or_tmp_111);
  assign and_131_cse = and_9_tmp & (fsm_output[1]);
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_cse = core_wen & (~((~ and_5_tmp)
      | (fsm_output[0])));
  assign and_11_cse = (~ plm_outputs_rsc_rls_obj_bawt) & exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_3;
  assign and_10_cse = (~ plm_outputs_rsci_bawt) & CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_3;
  assign COMPUTE_LOOP_buf_acc_data_and_cse = core_wen & (~ or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_j_and_cse = core_wen & and_7_tmp;
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_6_cse = core_wen & (~ or_tmp_111);
  assign CONVOLUTION_LOOP_for_for_for_for_for_n_and_itm = core_wen & and_9_tmp;
  assign CONVOLUTION_LOOP_for_and_3_rgt = (~ or_tmp_46) & and_dcpl_73;
  assign CONVOLUTION_LOOP_for_and_4_rgt = or_tmp_46 & and_dcpl_73;
  assign and_89_m1c = or_tmp_46 & and_9_tmp;
  assign and_88_rgt = (~ or_tmp_46) & and_9_tmp;
  assign CONVOLUTION_LOOP_for_for_and_3_rgt = (~ mux_35_cse) & and_89_m1c;
  assign CONVOLUTION_LOOP_for_for_and_4_rgt = mux_35_cse & and_89_m1c;
  assign and_91_m1c = mux_35_cse & and_9_tmp;
  assign and_90_rgt = (~ mux_35_cse) & and_9_tmp;
  assign CONVOLUTION_LOOP_for_for_for_and_2588_rgt = (~ mux_tmp_17) & and_91_m1c;
  assign CONVOLUTION_LOOP_for_for_for_and_2589_rgt = mux_tmp_17 & and_91_m1c;
  assign CONVOLUTION_LOOP_for_for_for_y_and_rgt = (~ and_dcpl_84) & and_dcpl_57;
  assign CONVOLUTION_LOOP_for_for_for_y_and_1_rgt = and_dcpl_84 & and_dcpl_57;
  assign exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0 = MUX_s_1_2_2(exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1,
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_1, and_7_tmp);
  assign lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0 = MUX_s_1_2_2(lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1,
      (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_1), and_7_tmp);
  assign CONVOLUTION_LOOP_CONVOLUTION_LOOP_CONVOLUTION_LOOP_COMPUTE_LOOP_not_1_nl
      = ~ COMPUTE_LOOP_COMPUTE_LOOP_or_tmp;
  assign CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0 = MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_4_0,
      CONVOLUTION_LOOP_CONVOLUTION_LOOP_CONVOLUTION_LOOP_COMPUTE_LOOP_not_1_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1954_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0,
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1, and_dcpl_66);
  assign exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_mx0w0 = CONVOLUTION_LOOP_for_for_for_for_mux_1954_nl
      & (~(operator_8_false_6_acc_itm_3_1 & ((~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp
      & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)) | (operator_8_false_1_acc_tmp[8]))));
  assign CONVOLUTION_LOOP_mux_6_nl = MUX_s_1_2_2(or_113_cse, exit_CONVOLUTION_LOOP_lpi_1_dfm_1,
      nand_tmp_7);
  assign exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0 = CONVOLUTION_LOOP_mux_6_nl & exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3_mx0w0;
  assign COMPUTE_LOOP_COMPUTE_LOOP_or_tmp = exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1
      | exit_COMPUTE_LOOP_lpi_1_dfm_2 | exitL_exit_COMPUTE_LOOP_sva;
  assign COMPUTE_LOOP_if_COMPUTE_LOOP_if_nand_tmp = ~((COMPUTE_LOOP_b_4_0_lpi_1_dfm_3_0_1
      == (operator_8_false_8_acc_tmp[3:0])) & (operator_8_false_8_acc_tmp[7:4]==4'b0000));
  assign exit_COMPUTE_LOOP_sva_2_mx0w0 = ~(COMPUTE_LOOP_if_COMPUTE_LOOP_if_nand_tmp
      | (operator_8_false_8_acc_tmp[8]));
  assign conf_info_crt_lpi_1_dfm_231_224_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_231_224,
      (conf_info_rsci_idat_mxwt[63:56]), exitL_exit_COMPUTE_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_71_64_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_71_64,
      (conf_info_rsci_idat_mxwt[23:16]), exitL_exit_COMPUTE_LOOP_sva);
  assign CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_if_CONVOLUTION_LOOP_for_if_nor_cse
      = ~((~(CONVOLUTION_LOOP_for_if_equal_tmp & (operator_8_false_3_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_3_acc_tmp[8]));
  assign exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1_mx0w0 = (CONVOLUTION_LOOP_for_acc_tmp[5])
      | CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_if_CONVOLUTION_LOOP_for_if_nor_cse;
  assign CONVOLUTION_LOOP_for_for_if_or_cse = (~((CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6
      == (operator_8_false_5_acc_tmp[4:0])) & (operator_8_false_5_acc_tmp[7:5]==3'b000)))
      | (operator_8_false_5_acc_tmp[8]);
  assign exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0 = ~(operator_8_false_3_acc_itm_4_1
      & CONVOLUTION_LOOP_for_for_if_or_cse);
  assign nl_if_acc_nl = if_acc_4_cse_1 + (conf_info_rsci_idat_mxwt[55:48]) + 8'b00000001;
  assign if_acc_nl = nl_if_acc_nl[7:0];
  assign operator_42_true_and_nl = (else_acc_psp_sva_1[10]) & (else_acc_psp_sva_1[0]);
  assign nl_operator_43_true_acc_nl = (else_acc_psp_sva_1[8:1]) + conv_u2s_1_8(operator_42_true_and_nl)
      + 8'b00000001;
  assign operator_43_true_acc_nl = nl_operator_43_true_acc_nl[7:0];
  assign n_w_out_lpi_1_dfm_3 = MUX1HOT_v_8_3_2(n_w_out_lpi_1_dfm_1, if_acc_nl, operator_43_true_acc_nl,
      {(~ exitL_exit_COMPUTE_LOOP_sva) , COMPUTE_LOOP_asn_44 , COMPUTE_LOOP_asn_46});
  assign nl_if_acc_6_nl = if_acc_4_cse_1 + (conf_info_rsci_idat_mxwt[47:40]) + 8'b00000001;
  assign if_acc_6_nl = nl_if_acc_6_nl[7:0];
  assign operator_42_true_1_and_nl = (else_acc_2_psp_sva_1[10]) & (else_acc_2_psp_sva_1[0]);
  assign nl_operator_43_true_1_acc_nl = (else_acc_2_psp_sva_1[8:1]) + conv_u2s_1_8(operator_42_true_1_and_nl)
      + 8'b00000001;
  assign operator_43_true_1_acc_nl = nl_operator_43_true_1_acc_nl[7:0];
  assign n_h_out_lpi_1_dfm_3 = MUX1HOT_v_8_3_2(n_h_out_lpi_1_dfm_1, if_acc_6_nl,
      operator_43_true_1_acc_nl, {(~ exitL_exit_COMPUTE_LOOP_sva) , COMPUTE_LOOP_asn_44
      , COMPUTE_LOOP_asn_46});
  assign conf_info_crt_lpi_1_dfm_135_128_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_135_128,
      (conf_info_rsci_idat_mxwt[39:32]), exitL_exit_COMPUTE_LOOP_sva);
  assign exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0 = ~(operator_8_false_5_acc_itm_3_1
      & ((~(CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp))
      | (operator_8_false_1_acc_tmp[8])));
  assign COMPUTE_LOOP_mux_4_nl = MUX_s_1_2_2(exit_COMPUTE_LOOP_sva_2_mx0w0, exit_COMPUTE_LOOP_sva_2,
      mux_tmp_21);
  assign exit_COMPUTE_LOOP_lpi_1_dfm_2_mx0w0 = ((COMPUTE_LOOP_acc_tmp[4]) | COMPUTE_LOOP_mux_4_nl)
      & exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0;
  assign CONVOLUTION_LOOP_for_mux_1_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1_mx0w0,
      exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1, or_tmp_46);
  assign exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3_mx0w0 = CONVOLUTION_LOOP_for_mux_1_nl
      & exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3_mx0w0;
  assign CONVOLUTION_LOOP_for_for_mux_1_nl = MUX_s_1_2_2(exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0,
      exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1, mux_35_cse);
  assign exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3_mx0w0 = CONVOLUTION_LOOP_for_for_mux_1_nl
      & exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_2_CONVOLUTION_LOOP_for_for_for_if_2_nor_cse
      = ~((~((CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6 == (operator_8_false_4_acc_tmp[4:0]))
      & (operator_8_false_4_acc_tmp[7:5]==3'b000))) | (operator_8_false_4_acc_tmp[8]));
  assign exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0 = (CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_2_CONVOLUTION_LOOP_for_for_for_if_2_nor_cse
      | (~ operator_8_false_4_acc_itm_4)) & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_mx0w0;
  assign conf_info_crt_lpi_1_dfm_103_96_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_103_96,
      (conf_info_rsci_idat_mxwt[31:24]), exitL_exit_COMPUTE_LOOP_sva);
  assign CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0 = ~((~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[0])
      | CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl = ~(MUX_v_45_2_2((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[45:1]),
      45'b111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0 = ~(MUX_v_45_2_2(CONVOLUTION_LOOP_for_for_for_for_for_nor_2_nl,
      45'b111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0 = ~((~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[46])
      | CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1);
  assign conf_info_crt_lpi_1_dfm_7_0_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_7_0,
      (conf_info_rsci_idat_mxwt[7:0]), exitL_exit_COMPUTE_LOOP_sva);
  assign CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp = CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_4
      == (operator_8_false_1_acc_tmp[2:0]);
  assign exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0 = exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0
      | (~((~ exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2) & lfst_exit_CONVOLUTION_LOOP_for_for_1_lpi_1_dfm_1));
  assign CONVOLUTION_LOOP_if_CONVOLUTION_LOOP_if_nand_tmp = ~((CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_4_0_1
      == (operator_8_false_7_acc_tmp[4:0])) & (operator_8_false_7_acc_tmp[7:5]==3'b000));
  assign CONVOLUTION_LOOP_for_if_equal_tmp = CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0
      == (operator_8_false_3_acc_tmp[4:0]);
  assign nl_n_w_in_acc_nl = (conf_info_rsci_idat_mxwt[55:49]) + (pad_sva_1[6:0]);
  assign n_w_in_acc_nl = nl_n_w_in_acc_nl[6:0];
  assign n_w_in_acc_psp_lpi_1_dfm_mx0 = MUX_v_7_2_2(n_w_in_acc_psp_lpi_1_dfm, n_w_in_acc_nl,
      exitL_exit_COMPUTE_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_192_mx0 = MUX_s_1_2_2(conf_info_crt_lpi_1_dfm_192,
      (conf_info_rsci_idat_mxwt[48]), exitL_exit_COMPUTE_LOOP_sva);
  assign nl_n_h_in_acc_nl = (conf_info_rsci_idat_mxwt[47:41]) + (pad_sva_1[6:0]);
  assign n_h_in_acc_nl = nl_n_h_in_acc_nl[6:0];
  assign n_h_in_acc_psp_lpi_1_dfm_mx0 = MUX_v_7_2_2(n_h_in_acc_psp_lpi_1_dfm, n_h_in_acc_nl,
      exitL_exit_COMPUTE_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_160_mx0 = MUX_s_1_2_2(conf_info_crt_lpi_1_dfm_160,
      (conf_info_rsci_idat_mxwt[40]), exitL_exit_COMPUTE_LOOP_sva);
  assign CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b00);
  assign CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[4:3]==2'b01);
  assign CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1 = ~((~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[0])
      | CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1)) | CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_nor_1_nl = ~(MUX_v_55_2_2((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[55:1]),
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0 = ~(MUX_v_55_2_2(CONVOLUTION_LOOP_for_for_for_else_nor_1_nl,
      55'b1111111111111111111111111111111111111111111111111111111, CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_67_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_66_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_65_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_64_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_63_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_62_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_61_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_60_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_59_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_58_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_57_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_56_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_55_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_54_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_53_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_52_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_51_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_50_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_49_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_48_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_47_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_46_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_45_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_44_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_43_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_42_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_41_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_40_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_7_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[3]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_127_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_68_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_126_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_69_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_125_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_70_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_124_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_71_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_123_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_72_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_122_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_73_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_121_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_74_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_120_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_75_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_119_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_76_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_118_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_77_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_117_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_78_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_116_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_79_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_115_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_80_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_114_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_81_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_113_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_82_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_112_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_83_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_111_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_84_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_110_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_85_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_109_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_86_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_108_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_87_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_107_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_88_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_106_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_89_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_105_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_90_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_104_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_91_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_103_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_92_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_102_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_93_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_101_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_94_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_100_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_95_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_99_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_96_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_98_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_97_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_67_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_66_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_65_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_64_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_63_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_62_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_61_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_60_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_59_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_58_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_57_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_56_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_55_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_54_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_53_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_52_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_51_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_50_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_49_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_48_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_47_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_46_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_45_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_44_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_43_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_42_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_41_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_40_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_6_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_32_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_33_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_34_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_35_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_36_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_37_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_38_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_39_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_40_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_41_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_42_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_43_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_44_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_45_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_46_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_47_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_48_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_49_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_50_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_51_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_52_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_53_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_54_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_55_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_56_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_57_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_58_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_59_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_60_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_61_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_62_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_63_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_5_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_16_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_17_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_18_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_19_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_20_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_21_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_22_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_23_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_24_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_25_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_26_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_27_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_28_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_29_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_30_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_31_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_4_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_8_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_9_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_10_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_11_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_12_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_13_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_14_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_15_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_3_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[2]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_4_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_5_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_6_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_7_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_0_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_1_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_2_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_2_3_sva_1 = CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[1]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_0_sva_1 = ~(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0
      | (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_1_sva_1 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0
      & (~ (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[0]));
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_2_sva_1 = (~ CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0)
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[0]);
  assign CONVOLUTION_LOOP_for_for_for_else_and_stg_1_3_sva_1 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0
      & (reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse[0]);
  assign nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1 = conv_s2s_57_58({CONVOLUTION_LOOP_for_for_for_else_mux_itm_1
      , CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1 , CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1})
      + conv_s2s_47_58({CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0 , CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0
      , CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0});
  assign CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:0];
  assign CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:56]==2'b10);
  assign CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[57:56]!=2'b01));
  assign CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_45_1_1
      = MUX_v_45_324_2(COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_3,
      {reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse , reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse
      , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0});
  assign CONVOLUTION_LOOP_for_for_for_if_1_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_56_46_1[10])
      & (~((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_45_1_1[44:30]==15'b111111111111111)
      & (CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_56_46_1[9:0]==10'b1111111111)));
  assign CONVOLUTION_LOOP_for_for_for_if_1_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_56_46_1[10])
      | (~((CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_45_1_1[44:30]!=15'b000000000000000)
      | (CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_56_46_1[9:0]!=10'b0000000000))));
  assign CONVOLUTION_LOOP_for_for_for_if_mux_974_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_978_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_974_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_978_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_975_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_980_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_975_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_980_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_976_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_982_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_976_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_982_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_977_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_984_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_977_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_984_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_978_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_986_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_978_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_986_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_979_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_988_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_979_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_988_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_980_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_990_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_980_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_990_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_981_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_992_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_981_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_992_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_982_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_994_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_982_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_994_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_983_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_996_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_983_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_996_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_984_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_998_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_984_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_998_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_985_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_985_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1000_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_986_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_986_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1002_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_987_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_987_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1004_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_988_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_988_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1006_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_989_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_989_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1008_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_990_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_990_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1010_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_991_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_991_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1012_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_992_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_992_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1014_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_993_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_993_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1016_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_994_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_994_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1018_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_995_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_995_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1020_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_996_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_996_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1022_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_997_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_997_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1024_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_998_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_998_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1026_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_999_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_999_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1028_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1000_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1030_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1001_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1032_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1002_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1034_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1003_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1036_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1004_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1038_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1005_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1040_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1006_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1042_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1007_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1044_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1008_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1046_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1009_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1048_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1010_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1050_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1011_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1052_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1012_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1054_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1013_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1056_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1014_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1058_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1015_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1060_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1016_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1062_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1017_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1064_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1018_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1066_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1019_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1068_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1020_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1070_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1021_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1072_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1022_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1074_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1023_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1076_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1024_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1078_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1025_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1080_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1026_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1082_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1027_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1084_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1028_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1086_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1029_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1088_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1030_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1090_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1031_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1092_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1032_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1094_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1033_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1096_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1034_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1098_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1035_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1100_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1036_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1102_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1037_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1104_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1038_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1106_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1039_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1108_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1040_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1110_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1041_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1112_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1042_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1114_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1043_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1116_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1044_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1118_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1045_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1120_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1046_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1122_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1047_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1124_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1048_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1126_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1049_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1128_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1050_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1130_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1051_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1132_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1052_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1134_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1053_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1136_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1054_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1138_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1055_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1140_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1056_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1142_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1057_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1144_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1058_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1146_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1059_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1148_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1060_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1150_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1061_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1152_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1062_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1154_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1063_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1156_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1064_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1158_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1065_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1160_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1066_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1162_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1067_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1164_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1068_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1166_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1069_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1168_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1070_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1170_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1071_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1172_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1072_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1174_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1073_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1176_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1074_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1178_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1075_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1180_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1076_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1182_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1077_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1184_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1078_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1186_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1079_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1188_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1080_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1190_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1081_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1192_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1082_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1194_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1083_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1196_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1084_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1198_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1085_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1200_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1086_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1202_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1087_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1204_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1088_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1206_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1089_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1208_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1090_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1210_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1091_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1212_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1092_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1214_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1093_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1216_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1094_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1218_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1095_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1220_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1096_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1222_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1097_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1224_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1098_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1226_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1099_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1228_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1100_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1230_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1101_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1232_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1102_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1234_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1103_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1236_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1104_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1238_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1105_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1240_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1106_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1242_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1107_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1244_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1108_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1246_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1109_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1248_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1110_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1250_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1111_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1252_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1112_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1254_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1113_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1256_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1114_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1258_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1115_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1260_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1116_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1262_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1117_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1264_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1118_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1266_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1119_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1268_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1120_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1270_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1121_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1272_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1122_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1274_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1123_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1276_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1124_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1278_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1125_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1280_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1126_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1282_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1127_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1284_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1128_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1286_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1129_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1288_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1130_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1290_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1131_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1292_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1132_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1294_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1133_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1296_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1134_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1298_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1135_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1300_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1136_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1302_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1137_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1304_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1138_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1306_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1139_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1308_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1140_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1310_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1141_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1312_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1142_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1314_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1143_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1316_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1144_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1318_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1145_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1320_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1146_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1322_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1147_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1324_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1148_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1326_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1149_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1328_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1150_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1330_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1151_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1332_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1152_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1334_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1153_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1336_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1154_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1338_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1155_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1340_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1156_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1342_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1157_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1344_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1158_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1346_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1159_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1348_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1160_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1350_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1161_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1352_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1162_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1354_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1163_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1356_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1164_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1358_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1165_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1360_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1166_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1362_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1167_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1364_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1168_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1366_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1169_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1368_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1170_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1370_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1171_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1372_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1172_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1374_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1173_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1376_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1174_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1378_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1175_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1380_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1176_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1382_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1177_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1384_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1178_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1386_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1179_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1388_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1180_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1390_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1181_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1392_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1182_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1394_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1183_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1396_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1184_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1398_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1185_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1400_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1186_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1402_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1187_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1404_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1188_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1406_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1189_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1408_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1190_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1410_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1191_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1412_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1192_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1414_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1193_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1416_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1194_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1418_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1195_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1420_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1196_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1422_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1197_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1424_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1198_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1426_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1199_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1428_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1200_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1430_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1201_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1432_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1202_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1434_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1203_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1436_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1204_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1438_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1205_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1440_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1206_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1442_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1207_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1444_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1208_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1446_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1209_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1448_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1210_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1450_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1211_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1452_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1212_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1454_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1213_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1456_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1214_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1458_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1215_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1460_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1216_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1462_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1217_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1464_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1218_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1466_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1219_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1468_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1220_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1470_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1221_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1472_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1222_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1474_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1223_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1476_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1224_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1478_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1225_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1480_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1226_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1482_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1227_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1484_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1228_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1486_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1229_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1488_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1230_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1490_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1231_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1492_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1232_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1494_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1233_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1496_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1234_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1498_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1235_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1500_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1236_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1502_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1237_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1504_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1238_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1506_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1239_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1508_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1240_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1510_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1241_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1512_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1242_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1514_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1243_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1516_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1244_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1518_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1245_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1520_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1246_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1522_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1247_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1524_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1248_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1526_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1249_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1528_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1250_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1530_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1251_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1532_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1252_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1534_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1253_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1536_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1254_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1538_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1255_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1540_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1256_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1542_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1257_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1544_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1258_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1546_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1259_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1548_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1260_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1550_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1261_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1552_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1262_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1554_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1263_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1556_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1264_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1558_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1265_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1560_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1266_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1562_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1267_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1564_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1268_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1566_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1269_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1568_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1270_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1570_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1271_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1572_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1272_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1574_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1273_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1576_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1274_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1578_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1275_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1580_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1276_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1582_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1277_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1584_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1278_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1586_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1279_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1588_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1280_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1590_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1281_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1592_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1282_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1594_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1283_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1596_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1284_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1598_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1285_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1600_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1286_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1602_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1287_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1604_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1288_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1606_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1289_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1608_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1290_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1610_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1291_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1612_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1292_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1614_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1293_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1616_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1294_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1618_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1295_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1620_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1296_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1622_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_mux_1297_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_0_sva_1, CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1);
  assign COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_if_mux_1297_nl,
      CONVOLUTION_LOOP_for_for_for_else_mux_1624_nl, CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_if_1_slc_COMPUTE_LOOP_buf_acc_data_57_56_0_sat_sva_56_46_1
      = MUX_v_11_324_2(COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_3, COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_3,
      {reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse , reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse
      , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0});
  assign COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5513
      , CONVOLUTION_LOOP_for_for_for_asn_5515 , CONVOLUTION_LOOP_for_for_for_asn_5517});
  assign COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5507
      , CONVOLUTION_LOOP_for_for_for_asn_5509 , CONVOLUTION_LOOP_for_for_for_asn_5511});
  assign COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5501
      , CONVOLUTION_LOOP_for_for_for_asn_5503 , CONVOLUTION_LOOP_for_for_for_asn_5505});
  assign COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5495
      , CONVOLUTION_LOOP_for_for_for_asn_5497 , CONVOLUTION_LOOP_for_for_for_asn_5499});
  assign COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5489
      , CONVOLUTION_LOOP_for_for_for_asn_5491 , CONVOLUTION_LOOP_for_for_for_asn_5493});
  assign COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5483
      , CONVOLUTION_LOOP_for_for_for_asn_5485 , CONVOLUTION_LOOP_for_for_for_asn_5487});
  assign COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5477
      , CONVOLUTION_LOOP_for_for_for_asn_5479 , CONVOLUTION_LOOP_for_for_for_asn_5481});
  assign COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5471
      , CONVOLUTION_LOOP_for_for_for_asn_5473 , CONVOLUTION_LOOP_for_for_for_asn_5475});
  assign COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5465
      , CONVOLUTION_LOOP_for_for_for_asn_5467 , CONVOLUTION_LOOP_for_for_for_asn_5469});
  assign COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5459
      , CONVOLUTION_LOOP_for_for_for_asn_5461 , CONVOLUTION_LOOP_for_for_for_asn_5463});
  assign COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5453
      , CONVOLUTION_LOOP_for_for_for_asn_5455 , CONVOLUTION_LOOP_for_for_for_asn_5457});
  assign COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5447
      , CONVOLUTION_LOOP_for_for_for_asn_5449 , CONVOLUTION_LOOP_for_for_for_asn_5451});
  assign COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5441
      , CONVOLUTION_LOOP_for_for_for_asn_5443 , CONVOLUTION_LOOP_for_for_for_asn_5445});
  assign COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5435
      , CONVOLUTION_LOOP_for_for_for_asn_5437 , CONVOLUTION_LOOP_for_for_for_asn_5439});
  assign COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5429
      , CONVOLUTION_LOOP_for_for_for_asn_5431 , CONVOLUTION_LOOP_for_for_for_asn_5433});
  assign COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5423
      , CONVOLUTION_LOOP_for_for_for_asn_5425 , CONVOLUTION_LOOP_for_for_for_asn_5427});
  assign COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5417
      , CONVOLUTION_LOOP_for_for_for_asn_5419 , CONVOLUTION_LOOP_for_for_for_asn_5421});
  assign COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5411
      , CONVOLUTION_LOOP_for_for_for_asn_5413 , CONVOLUTION_LOOP_for_for_for_asn_5415});
  assign COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5405
      , CONVOLUTION_LOOP_for_for_for_asn_5407 , CONVOLUTION_LOOP_for_for_for_asn_5409});
  assign COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5399
      , CONVOLUTION_LOOP_for_for_for_asn_5401 , CONVOLUTION_LOOP_for_for_for_asn_5403});
  assign COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5393
      , CONVOLUTION_LOOP_for_for_for_asn_5395 , CONVOLUTION_LOOP_for_for_for_asn_5397});
  assign COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5387
      , CONVOLUTION_LOOP_for_for_for_asn_5389 , CONVOLUTION_LOOP_for_for_for_asn_5391});
  assign COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5381
      , CONVOLUTION_LOOP_for_for_for_asn_5383 , CONVOLUTION_LOOP_for_for_for_asn_5385});
  assign COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5375
      , CONVOLUTION_LOOP_for_for_for_asn_5377 , CONVOLUTION_LOOP_for_for_for_asn_5379});
  assign COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5369
      , CONVOLUTION_LOOP_for_for_for_asn_5371 , CONVOLUTION_LOOP_for_for_for_asn_5373});
  assign COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5363
      , CONVOLUTION_LOOP_for_for_for_asn_5365 , CONVOLUTION_LOOP_for_for_for_asn_5367});
  assign COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5357
      , CONVOLUTION_LOOP_for_for_for_asn_5359 , CONVOLUTION_LOOP_for_for_for_asn_5361});
  assign COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5351
      , CONVOLUTION_LOOP_for_for_for_asn_5353 , CONVOLUTION_LOOP_for_for_for_asn_5355});
  assign COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5345
      , CONVOLUTION_LOOP_for_for_for_asn_5347 , CONVOLUTION_LOOP_for_for_for_asn_5349});
  assign COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5339
      , CONVOLUTION_LOOP_for_for_for_asn_5341 , CONVOLUTION_LOOP_for_for_for_asn_5343});
  assign COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5333
      , CONVOLUTION_LOOP_for_for_for_asn_5335 , CONVOLUTION_LOOP_for_for_for_asn_5337});
  assign COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5327
      , CONVOLUTION_LOOP_for_for_for_asn_5329 , CONVOLUTION_LOOP_for_for_for_asn_5331});
  assign COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5321
      , CONVOLUTION_LOOP_for_for_for_asn_5323 , CONVOLUTION_LOOP_for_for_for_asn_5325});
  assign COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5315
      , CONVOLUTION_LOOP_for_for_for_asn_5317 , CONVOLUTION_LOOP_for_for_for_asn_5319});
  assign COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5309
      , CONVOLUTION_LOOP_for_for_for_asn_5311 , CONVOLUTION_LOOP_for_for_for_asn_5313});
  assign COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5303
      , CONVOLUTION_LOOP_for_for_for_asn_5305 , CONVOLUTION_LOOP_for_for_for_asn_5307});
  assign COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5297
      , CONVOLUTION_LOOP_for_for_for_asn_5299 , CONVOLUTION_LOOP_for_for_for_asn_5301});
  assign COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5291
      , CONVOLUTION_LOOP_for_for_for_asn_5293 , CONVOLUTION_LOOP_for_for_for_asn_5295});
  assign COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5285
      , CONVOLUTION_LOOP_for_for_for_asn_5287 , CONVOLUTION_LOOP_for_for_for_asn_5289});
  assign COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5279
      , CONVOLUTION_LOOP_for_for_for_asn_5281 , CONVOLUTION_LOOP_for_for_for_asn_5283});
  assign COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5273
      , CONVOLUTION_LOOP_for_for_for_asn_5275 , CONVOLUTION_LOOP_for_for_for_asn_5277});
  assign COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5267
      , CONVOLUTION_LOOP_for_for_for_asn_5269 , CONVOLUTION_LOOP_for_for_for_asn_5271});
  assign COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5261
      , CONVOLUTION_LOOP_for_for_for_asn_5263 , CONVOLUTION_LOOP_for_for_for_asn_5265});
  assign COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5255
      , CONVOLUTION_LOOP_for_for_for_asn_5257 , CONVOLUTION_LOOP_for_for_for_asn_5259});
  assign COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5249
      , CONVOLUTION_LOOP_for_for_for_asn_5251 , CONVOLUTION_LOOP_for_for_for_asn_5253});
  assign COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5243
      , CONVOLUTION_LOOP_for_for_for_asn_5245 , CONVOLUTION_LOOP_for_for_for_asn_5247});
  assign COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5237
      , CONVOLUTION_LOOP_for_for_for_asn_5239 , CONVOLUTION_LOOP_for_for_for_asn_5241});
  assign COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5231
      , CONVOLUTION_LOOP_for_for_for_asn_5233 , CONVOLUTION_LOOP_for_for_for_asn_5235});
  assign COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5225
      , CONVOLUTION_LOOP_for_for_for_asn_5227 , CONVOLUTION_LOOP_for_for_for_asn_5229});
  assign COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5219
      , CONVOLUTION_LOOP_for_for_for_asn_5221 , CONVOLUTION_LOOP_for_for_for_asn_5223});
  assign COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5213
      , CONVOLUTION_LOOP_for_for_for_asn_5215 , CONVOLUTION_LOOP_for_for_for_asn_5217});
  assign COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5207
      , CONVOLUTION_LOOP_for_for_for_asn_5209 , CONVOLUTION_LOOP_for_for_for_asn_5211});
  assign COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5201
      , CONVOLUTION_LOOP_for_for_for_asn_5203 , CONVOLUTION_LOOP_for_for_for_asn_5205});
  assign COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5195
      , CONVOLUTION_LOOP_for_for_for_asn_5197 , CONVOLUTION_LOOP_for_for_for_asn_5199});
  assign COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5189
      , CONVOLUTION_LOOP_for_for_for_asn_5191 , CONVOLUTION_LOOP_for_for_for_asn_5193});
  assign COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5183
      , CONVOLUTION_LOOP_for_for_for_asn_5185 , CONVOLUTION_LOOP_for_for_for_asn_5187});
  assign COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5177
      , CONVOLUTION_LOOP_for_for_for_asn_5179 , CONVOLUTION_LOOP_for_for_for_asn_5181});
  assign COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5171
      , CONVOLUTION_LOOP_for_for_for_asn_5173 , CONVOLUTION_LOOP_for_for_for_asn_5175});
  assign COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5165
      , CONVOLUTION_LOOP_for_for_for_asn_5167 , CONVOLUTION_LOOP_for_for_for_asn_5169});
  assign COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5159
      , CONVOLUTION_LOOP_for_for_for_asn_5161 , CONVOLUTION_LOOP_for_for_for_asn_5163});
  assign COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5153
      , CONVOLUTION_LOOP_for_for_for_asn_5155 , CONVOLUTION_LOOP_for_for_for_asn_5157});
  assign COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5147
      , CONVOLUTION_LOOP_for_for_for_asn_5149 , CONVOLUTION_LOOP_for_for_for_asn_5151});
  assign COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5141
      , CONVOLUTION_LOOP_for_for_for_asn_5143 , CONVOLUTION_LOOP_for_for_for_asn_5145});
  assign COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5135
      , CONVOLUTION_LOOP_for_for_for_asn_5137 , CONVOLUTION_LOOP_for_for_for_asn_5139});
  assign COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5129
      , CONVOLUTION_LOOP_for_for_for_asn_5131 , CONVOLUTION_LOOP_for_for_for_asn_5133});
  assign COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5123
      , CONVOLUTION_LOOP_for_for_for_asn_5125 , CONVOLUTION_LOOP_for_for_for_asn_5127});
  assign COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5117
      , CONVOLUTION_LOOP_for_for_for_asn_5119 , CONVOLUTION_LOOP_for_for_for_asn_5121});
  assign COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5111
      , CONVOLUTION_LOOP_for_for_for_asn_5113 , CONVOLUTION_LOOP_for_for_for_asn_5115});
  assign COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5105
      , CONVOLUTION_LOOP_for_for_for_asn_5107 , CONVOLUTION_LOOP_for_for_for_asn_5109});
  assign COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5099
      , CONVOLUTION_LOOP_for_for_for_asn_5101 , CONVOLUTION_LOOP_for_for_for_asn_5103});
  assign COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5093
      , CONVOLUTION_LOOP_for_for_for_asn_5095 , CONVOLUTION_LOOP_for_for_for_asn_5097});
  assign COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5087
      , CONVOLUTION_LOOP_for_for_for_asn_5089 , CONVOLUTION_LOOP_for_for_for_asn_5091});
  assign COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5081
      , CONVOLUTION_LOOP_for_for_for_asn_5083 , CONVOLUTION_LOOP_for_for_for_asn_5085});
  assign COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5075
      , CONVOLUTION_LOOP_for_for_for_asn_5077 , CONVOLUTION_LOOP_for_for_for_asn_5079});
  assign COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5069
      , CONVOLUTION_LOOP_for_for_for_asn_5071 , CONVOLUTION_LOOP_for_for_for_asn_5073});
  assign COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5063
      , CONVOLUTION_LOOP_for_for_for_asn_5065 , CONVOLUTION_LOOP_for_for_for_asn_5067});
  assign COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5057
      , CONVOLUTION_LOOP_for_for_for_asn_5059 , CONVOLUTION_LOOP_for_for_for_asn_5061});
  assign COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5051
      , CONVOLUTION_LOOP_for_for_for_asn_5053 , CONVOLUTION_LOOP_for_for_for_asn_5055});
  assign COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5045
      , CONVOLUTION_LOOP_for_for_for_asn_5047 , CONVOLUTION_LOOP_for_for_for_asn_5049});
  assign COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5039
      , CONVOLUTION_LOOP_for_for_for_asn_5041 , CONVOLUTION_LOOP_for_for_for_asn_5043});
  assign COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5033
      , CONVOLUTION_LOOP_for_for_for_asn_5035 , CONVOLUTION_LOOP_for_for_for_asn_5037});
  assign COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5027
      , CONVOLUTION_LOOP_for_for_for_asn_5029 , CONVOLUTION_LOOP_for_for_for_asn_5031});
  assign COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5021
      , CONVOLUTION_LOOP_for_for_for_asn_5023 , CONVOLUTION_LOOP_for_for_for_asn_5025});
  assign COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5015
      , CONVOLUTION_LOOP_for_for_for_asn_5017 , CONVOLUTION_LOOP_for_for_for_asn_5019});
  assign COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5009
      , CONVOLUTION_LOOP_for_for_for_asn_5011 , CONVOLUTION_LOOP_for_for_for_asn_5013});
  assign COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_5003
      , CONVOLUTION_LOOP_for_for_for_asn_5005 , CONVOLUTION_LOOP_for_for_for_asn_5007});
  assign COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4997
      , CONVOLUTION_LOOP_for_for_for_asn_4999 , CONVOLUTION_LOOP_for_for_for_asn_5001});
  assign COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4991
      , CONVOLUTION_LOOP_for_for_for_asn_4993 , CONVOLUTION_LOOP_for_for_for_asn_4995});
  assign COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4985
      , CONVOLUTION_LOOP_for_for_for_asn_4987 , CONVOLUTION_LOOP_for_for_for_asn_4989});
  assign COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4979
      , CONVOLUTION_LOOP_for_for_for_asn_4981 , CONVOLUTION_LOOP_for_for_for_asn_4983});
  assign COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4973
      , CONVOLUTION_LOOP_for_for_for_asn_4975 , CONVOLUTION_LOOP_for_for_for_asn_4977});
  assign COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4967
      , CONVOLUTION_LOOP_for_for_for_asn_4969 , CONVOLUTION_LOOP_for_for_for_asn_4971});
  assign COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4961
      , CONVOLUTION_LOOP_for_for_for_asn_4963 , CONVOLUTION_LOOP_for_for_for_asn_4965});
  assign COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4955
      , CONVOLUTION_LOOP_for_for_for_asn_4957 , CONVOLUTION_LOOP_for_for_for_asn_4959});
  assign COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4949
      , CONVOLUTION_LOOP_for_for_for_asn_4951 , CONVOLUTION_LOOP_for_for_for_asn_4953});
  assign COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4943
      , CONVOLUTION_LOOP_for_for_for_asn_4945 , CONVOLUTION_LOOP_for_for_for_asn_4947});
  assign COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4937
      , CONVOLUTION_LOOP_for_for_for_asn_4939 , CONVOLUTION_LOOP_for_for_for_asn_4941});
  assign COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4931
      , CONVOLUTION_LOOP_for_for_for_asn_4933 , CONVOLUTION_LOOP_for_for_for_asn_4935});
  assign COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4925
      , CONVOLUTION_LOOP_for_for_for_asn_4927 , CONVOLUTION_LOOP_for_for_for_asn_4929});
  assign COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4919
      , CONVOLUTION_LOOP_for_for_for_asn_4921 , CONVOLUTION_LOOP_for_for_for_asn_4923});
  assign COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4913
      , CONVOLUTION_LOOP_for_for_for_asn_4915 , CONVOLUTION_LOOP_for_for_for_asn_4917});
  assign COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4907
      , CONVOLUTION_LOOP_for_for_for_asn_4909 , CONVOLUTION_LOOP_for_for_for_asn_4911});
  assign COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4901
      , CONVOLUTION_LOOP_for_for_for_asn_4903 , CONVOLUTION_LOOP_for_for_for_asn_4905});
  assign COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4895
      , CONVOLUTION_LOOP_for_for_for_asn_4897 , CONVOLUTION_LOOP_for_for_for_asn_4899});
  assign COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4889
      , CONVOLUTION_LOOP_for_for_for_asn_4891 , CONVOLUTION_LOOP_for_for_for_asn_4893});
  assign COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4883
      , CONVOLUTION_LOOP_for_for_for_asn_4885 , CONVOLUTION_LOOP_for_for_for_asn_4887});
  assign COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4877
      , CONVOLUTION_LOOP_for_for_for_asn_4879 , CONVOLUTION_LOOP_for_for_for_asn_4881});
  assign COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4871
      , CONVOLUTION_LOOP_for_for_for_asn_4873 , CONVOLUTION_LOOP_for_for_for_asn_4875});
  assign COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4865
      , CONVOLUTION_LOOP_for_for_for_asn_4867 , CONVOLUTION_LOOP_for_for_for_asn_4869});
  assign COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4859
      , CONVOLUTION_LOOP_for_for_for_asn_4861 , CONVOLUTION_LOOP_for_for_for_asn_4863});
  assign COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4853
      , CONVOLUTION_LOOP_for_for_for_asn_4855 , CONVOLUTION_LOOP_for_for_for_asn_4857});
  assign COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4847
      , CONVOLUTION_LOOP_for_for_for_asn_4849 , CONVOLUTION_LOOP_for_for_for_asn_4851});
  assign COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4841
      , CONVOLUTION_LOOP_for_for_for_asn_4843 , CONVOLUTION_LOOP_for_for_for_asn_4845});
  assign COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4835
      , CONVOLUTION_LOOP_for_for_for_asn_4837 , CONVOLUTION_LOOP_for_for_for_asn_4839});
  assign COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4829
      , CONVOLUTION_LOOP_for_for_for_asn_4831 , CONVOLUTION_LOOP_for_for_for_asn_4833});
  assign COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4823
      , CONVOLUTION_LOOP_for_for_for_asn_4825 , CONVOLUTION_LOOP_for_for_for_asn_4827});
  assign COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4817
      , CONVOLUTION_LOOP_for_for_for_asn_4819 , CONVOLUTION_LOOP_for_for_for_asn_4821});
  assign COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4811
      , CONVOLUTION_LOOP_for_for_for_asn_4813 , CONVOLUTION_LOOP_for_for_for_asn_4815});
  assign COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4805
      , CONVOLUTION_LOOP_for_for_for_asn_4807 , CONVOLUTION_LOOP_for_for_for_asn_4809});
  assign COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4799
      , CONVOLUTION_LOOP_for_for_for_asn_4801 , CONVOLUTION_LOOP_for_for_for_asn_4803});
  assign COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4793
      , CONVOLUTION_LOOP_for_for_for_asn_4795 , CONVOLUTION_LOOP_for_for_for_asn_4797});
  assign COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4787
      , CONVOLUTION_LOOP_for_for_for_asn_4789 , CONVOLUTION_LOOP_for_for_for_asn_4791});
  assign COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4781
      , CONVOLUTION_LOOP_for_for_for_asn_4783 , CONVOLUTION_LOOP_for_for_for_asn_4785});
  assign COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4775
      , CONVOLUTION_LOOP_for_for_for_asn_4777 , CONVOLUTION_LOOP_for_for_for_asn_4779});
  assign COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4769
      , CONVOLUTION_LOOP_for_for_for_asn_4771 , CONVOLUTION_LOOP_for_for_for_asn_4773});
  assign COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4763
      , CONVOLUTION_LOOP_for_for_for_asn_4765 , CONVOLUTION_LOOP_for_for_for_asn_4767});
  assign COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4757
      , CONVOLUTION_LOOP_for_for_for_asn_4759 , CONVOLUTION_LOOP_for_for_for_asn_4761});
  assign COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4751
      , CONVOLUTION_LOOP_for_for_for_asn_4753 , CONVOLUTION_LOOP_for_for_for_asn_4755});
  assign COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4745
      , CONVOLUTION_LOOP_for_for_for_asn_4747 , CONVOLUTION_LOOP_for_for_for_asn_4749});
  assign COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4739
      , CONVOLUTION_LOOP_for_for_for_asn_4741 , CONVOLUTION_LOOP_for_for_for_asn_4743});
  assign COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4733
      , CONVOLUTION_LOOP_for_for_for_asn_4735 , CONVOLUTION_LOOP_for_for_for_asn_4737});
  assign COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4727
      , CONVOLUTION_LOOP_for_for_for_asn_4729 , CONVOLUTION_LOOP_for_for_for_asn_4731});
  assign COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4721
      , CONVOLUTION_LOOP_for_for_for_asn_4723 , CONVOLUTION_LOOP_for_for_for_asn_4725});
  assign COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4715
      , CONVOLUTION_LOOP_for_for_for_asn_4717 , CONVOLUTION_LOOP_for_for_for_asn_4719});
  assign COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4709
      , CONVOLUTION_LOOP_for_for_for_asn_4711 , CONVOLUTION_LOOP_for_for_for_asn_4713});
  assign COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4703
      , CONVOLUTION_LOOP_for_for_for_asn_4705 , CONVOLUTION_LOOP_for_for_for_asn_4707});
  assign COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4697
      , CONVOLUTION_LOOP_for_for_for_asn_4699 , CONVOLUTION_LOOP_for_for_for_asn_4701});
  assign COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4691
      , CONVOLUTION_LOOP_for_for_for_asn_4693 , CONVOLUTION_LOOP_for_for_for_asn_4695});
  assign COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4685
      , CONVOLUTION_LOOP_for_for_for_asn_4687 , CONVOLUTION_LOOP_for_for_for_asn_4689});
  assign COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4679
      , CONVOLUTION_LOOP_for_for_for_asn_4681 , CONVOLUTION_LOOP_for_for_for_asn_4683});
  assign COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4673
      , CONVOLUTION_LOOP_for_for_for_asn_4675 , CONVOLUTION_LOOP_for_for_for_asn_4677});
  assign COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4667
      , CONVOLUTION_LOOP_for_for_for_asn_4669 , CONVOLUTION_LOOP_for_for_for_asn_4671});
  assign COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4661
      , CONVOLUTION_LOOP_for_for_for_asn_4663 , CONVOLUTION_LOOP_for_for_for_asn_4665});
  assign COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4655
      , CONVOLUTION_LOOP_for_for_for_asn_4657 , CONVOLUTION_LOOP_for_for_for_asn_4659});
  assign COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4649
      , CONVOLUTION_LOOP_for_for_for_asn_4651 , CONVOLUTION_LOOP_for_for_for_asn_4653});
  assign COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4643
      , CONVOLUTION_LOOP_for_for_for_asn_4645 , CONVOLUTION_LOOP_for_for_for_asn_4647});
  assign COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4637
      , CONVOLUTION_LOOP_for_for_for_asn_4639 , CONVOLUTION_LOOP_for_for_for_asn_4641});
  assign COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4631
      , CONVOLUTION_LOOP_for_for_for_asn_4633 , CONVOLUTION_LOOP_for_for_for_asn_4635});
  assign COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4625
      , CONVOLUTION_LOOP_for_for_for_asn_4627 , CONVOLUTION_LOOP_for_for_for_asn_4629});
  assign COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4619
      , CONVOLUTION_LOOP_for_for_for_asn_4621 , CONVOLUTION_LOOP_for_for_for_asn_4623});
  assign COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4613
      , CONVOLUTION_LOOP_for_for_for_asn_4615 , CONVOLUTION_LOOP_for_for_for_asn_4617});
  assign COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4607
      , CONVOLUTION_LOOP_for_for_for_asn_4609 , CONVOLUTION_LOOP_for_for_for_asn_4611});
  assign COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4601
      , CONVOLUTION_LOOP_for_for_for_asn_4603 , CONVOLUTION_LOOP_for_for_for_asn_4605});
  assign COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4595
      , CONVOLUTION_LOOP_for_for_for_asn_4597 , CONVOLUTION_LOOP_for_for_for_asn_4599});
  assign COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4589
      , CONVOLUTION_LOOP_for_for_for_asn_4591 , CONVOLUTION_LOOP_for_for_for_asn_4593});
  assign COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4583
      , CONVOLUTION_LOOP_for_for_for_asn_4585 , CONVOLUTION_LOOP_for_for_for_asn_4587});
  assign COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4577
      , CONVOLUTION_LOOP_for_for_for_asn_4579 , CONVOLUTION_LOOP_for_for_for_asn_4581});
  assign COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4571
      , CONVOLUTION_LOOP_for_for_for_asn_4573 , CONVOLUTION_LOOP_for_for_for_asn_4575});
  assign COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4565
      , CONVOLUTION_LOOP_for_for_for_asn_4567 , CONVOLUTION_LOOP_for_for_for_asn_4569});
  assign COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4559
      , CONVOLUTION_LOOP_for_for_for_asn_4561 , CONVOLUTION_LOOP_for_for_for_asn_4563});
  assign COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4553
      , CONVOLUTION_LOOP_for_for_for_asn_4555 , CONVOLUTION_LOOP_for_for_for_asn_4557});
  assign COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4547
      , CONVOLUTION_LOOP_for_for_for_asn_4549 , CONVOLUTION_LOOP_for_for_for_asn_4551});
  assign COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4541
      , CONVOLUTION_LOOP_for_for_for_asn_4543 , CONVOLUTION_LOOP_for_for_for_asn_4545});
  assign COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4535
      , CONVOLUTION_LOOP_for_for_for_asn_4537 , CONVOLUTION_LOOP_for_for_for_asn_4539});
  assign COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4529
      , CONVOLUTION_LOOP_for_for_for_asn_4531 , CONVOLUTION_LOOP_for_for_for_asn_4533});
  assign COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4523
      , CONVOLUTION_LOOP_for_for_for_asn_4525 , CONVOLUTION_LOOP_for_for_for_asn_4527});
  assign COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4517
      , CONVOLUTION_LOOP_for_for_for_asn_4519 , CONVOLUTION_LOOP_for_for_for_asn_4521});
  assign COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4511
      , CONVOLUTION_LOOP_for_for_for_asn_4513 , CONVOLUTION_LOOP_for_for_for_asn_4515});
  assign COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4505
      , CONVOLUTION_LOOP_for_for_for_asn_4507 , CONVOLUTION_LOOP_for_for_for_asn_4509});
  assign COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4499
      , CONVOLUTION_LOOP_for_for_for_asn_4501 , CONVOLUTION_LOOP_for_for_for_asn_4503});
  assign COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4493
      , CONVOLUTION_LOOP_for_for_for_asn_4495 , CONVOLUTION_LOOP_for_for_for_asn_4497});
  assign COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4487
      , CONVOLUTION_LOOP_for_for_for_asn_4489 , CONVOLUTION_LOOP_for_for_for_asn_4491});
  assign COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4481
      , CONVOLUTION_LOOP_for_for_for_asn_4483 , CONVOLUTION_LOOP_for_for_for_asn_4485});
  assign COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4475
      , CONVOLUTION_LOOP_for_for_for_asn_4477 , CONVOLUTION_LOOP_for_for_for_asn_4479});
  assign COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4469
      , CONVOLUTION_LOOP_for_for_for_asn_4471 , CONVOLUTION_LOOP_for_for_for_asn_4473});
  assign COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4463
      , CONVOLUTION_LOOP_for_for_for_asn_4465 , CONVOLUTION_LOOP_for_for_for_asn_4467});
  assign COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4457
      , CONVOLUTION_LOOP_for_for_for_asn_4459 , CONVOLUTION_LOOP_for_for_for_asn_4461});
  assign COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4451
      , CONVOLUTION_LOOP_for_for_for_asn_4453 , CONVOLUTION_LOOP_for_for_for_asn_4455});
  assign COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4445
      , CONVOLUTION_LOOP_for_for_for_asn_4447 , CONVOLUTION_LOOP_for_for_for_asn_4449});
  assign COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4439
      , CONVOLUTION_LOOP_for_for_for_asn_4441 , CONVOLUTION_LOOP_for_for_for_asn_4443});
  assign COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4433
      , CONVOLUTION_LOOP_for_for_for_asn_4435 , CONVOLUTION_LOOP_for_for_for_asn_4437});
  assign COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4427
      , CONVOLUTION_LOOP_for_for_for_asn_4429 , CONVOLUTION_LOOP_for_for_for_asn_4431});
  assign COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4421
      , CONVOLUTION_LOOP_for_for_for_asn_4423 , CONVOLUTION_LOOP_for_for_for_asn_4425});
  assign COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4415
      , CONVOLUTION_LOOP_for_for_for_asn_4417 , CONVOLUTION_LOOP_for_for_for_asn_4419});
  assign COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4409
      , CONVOLUTION_LOOP_for_for_for_asn_4411 , CONVOLUTION_LOOP_for_for_for_asn_4413});
  assign COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4403
      , CONVOLUTION_LOOP_for_for_for_asn_4405 , CONVOLUTION_LOOP_for_for_for_asn_4407});
  assign COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4397
      , CONVOLUTION_LOOP_for_for_for_asn_4399 , CONVOLUTION_LOOP_for_for_for_asn_4401});
  assign COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4391
      , CONVOLUTION_LOOP_for_for_for_asn_4393 , CONVOLUTION_LOOP_for_for_for_asn_4395});
  assign COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4385
      , CONVOLUTION_LOOP_for_for_for_asn_4387 , CONVOLUTION_LOOP_for_for_for_asn_4389});
  assign COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4379
      , CONVOLUTION_LOOP_for_for_for_asn_4381 , CONVOLUTION_LOOP_for_for_for_asn_4383});
  assign COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4373
      , CONVOLUTION_LOOP_for_for_for_asn_4375 , CONVOLUTION_LOOP_for_for_for_asn_4377});
  assign COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4367
      , CONVOLUTION_LOOP_for_for_for_asn_4369 , CONVOLUTION_LOOP_for_for_for_asn_4371});
  assign COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4361
      , CONVOLUTION_LOOP_for_for_for_asn_4363 , CONVOLUTION_LOOP_for_for_for_asn_4365});
  assign COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4355
      , CONVOLUTION_LOOP_for_for_for_asn_4357 , CONVOLUTION_LOOP_for_for_for_asn_4359});
  assign COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4349
      , CONVOLUTION_LOOP_for_for_for_asn_4351 , CONVOLUTION_LOOP_for_for_for_asn_4353});
  assign COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4343
      , CONVOLUTION_LOOP_for_for_for_asn_4345 , CONVOLUTION_LOOP_for_for_for_asn_4347});
  assign COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4337
      , CONVOLUTION_LOOP_for_for_for_asn_4339 , CONVOLUTION_LOOP_for_for_for_asn_4341});
  assign COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4331
      , CONVOLUTION_LOOP_for_for_for_asn_4333 , CONVOLUTION_LOOP_for_for_for_asn_4335});
  assign COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4325
      , CONVOLUTION_LOOP_for_for_for_asn_4327 , CONVOLUTION_LOOP_for_for_for_asn_4329});
  assign COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4319
      , CONVOLUTION_LOOP_for_for_for_asn_4321 , CONVOLUTION_LOOP_for_for_for_asn_4323});
  assign COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4313
      , CONVOLUTION_LOOP_for_for_for_asn_4315 , CONVOLUTION_LOOP_for_for_for_asn_4317});
  assign COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4307
      , CONVOLUTION_LOOP_for_for_for_asn_4309 , CONVOLUTION_LOOP_for_for_for_asn_4311});
  assign COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4301
      , CONVOLUTION_LOOP_for_for_for_asn_4303 , CONVOLUTION_LOOP_for_for_for_asn_4305});
  assign COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4295
      , CONVOLUTION_LOOP_for_for_for_asn_4297 , CONVOLUTION_LOOP_for_for_for_asn_4299});
  assign COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4289
      , CONVOLUTION_LOOP_for_for_for_asn_4291 , CONVOLUTION_LOOP_for_for_for_asn_4293});
  assign COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4283
      , CONVOLUTION_LOOP_for_for_for_asn_4285 , CONVOLUTION_LOOP_for_for_for_asn_4287});
  assign COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4277
      , CONVOLUTION_LOOP_for_for_for_asn_4279 , CONVOLUTION_LOOP_for_for_for_asn_4281});
  assign COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4271
      , CONVOLUTION_LOOP_for_for_for_asn_4273 , CONVOLUTION_LOOP_for_for_for_asn_4275});
  assign COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4265
      , CONVOLUTION_LOOP_for_for_for_asn_4267 , CONVOLUTION_LOOP_for_for_for_asn_4269});
  assign COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4259
      , CONVOLUTION_LOOP_for_for_for_asn_4261 , CONVOLUTION_LOOP_for_for_for_asn_4263});
  assign COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4253
      , CONVOLUTION_LOOP_for_for_for_asn_4255 , CONVOLUTION_LOOP_for_for_for_asn_4257});
  assign COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4247
      , CONVOLUTION_LOOP_for_for_for_asn_4249 , CONVOLUTION_LOOP_for_for_for_asn_4251});
  assign COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4241
      , CONVOLUTION_LOOP_for_for_for_asn_4243 , CONVOLUTION_LOOP_for_for_for_asn_4245});
  assign COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4235
      , CONVOLUTION_LOOP_for_for_for_asn_4237 , CONVOLUTION_LOOP_for_for_for_asn_4239});
  assign COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4229
      , CONVOLUTION_LOOP_for_for_for_asn_4231 , CONVOLUTION_LOOP_for_for_for_asn_4233});
  assign COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4223
      , CONVOLUTION_LOOP_for_for_for_asn_4225 , CONVOLUTION_LOOP_for_for_for_asn_4227});
  assign COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4217
      , CONVOLUTION_LOOP_for_for_for_asn_4219 , CONVOLUTION_LOOP_for_for_for_asn_4221});
  assign COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4211
      , CONVOLUTION_LOOP_for_for_for_asn_4213 , CONVOLUTION_LOOP_for_for_for_asn_4215});
  assign COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4205
      , CONVOLUTION_LOOP_for_for_for_asn_4207 , CONVOLUTION_LOOP_for_for_for_asn_4209});
  assign COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4199
      , CONVOLUTION_LOOP_for_for_for_asn_4201 , CONVOLUTION_LOOP_for_for_for_asn_4203});
  assign COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4193
      , CONVOLUTION_LOOP_for_for_for_asn_4195 , CONVOLUTION_LOOP_for_for_for_asn_4197});
  assign COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4187
      , CONVOLUTION_LOOP_for_for_for_asn_4189 , CONVOLUTION_LOOP_for_for_for_asn_4191});
  assign COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4181
      , CONVOLUTION_LOOP_for_for_for_asn_4183 , CONVOLUTION_LOOP_for_for_for_asn_4185});
  assign COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4175
      , CONVOLUTION_LOOP_for_for_for_asn_4177 , CONVOLUTION_LOOP_for_for_for_asn_4179});
  assign COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4169
      , CONVOLUTION_LOOP_for_for_for_asn_4171 , CONVOLUTION_LOOP_for_for_for_asn_4173});
  assign COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4163
      , CONVOLUTION_LOOP_for_for_for_asn_4165 , CONVOLUTION_LOOP_for_for_for_asn_4167});
  assign COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4157
      , CONVOLUTION_LOOP_for_for_for_asn_4159 , CONVOLUTION_LOOP_for_for_for_asn_4161});
  assign COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4151
      , CONVOLUTION_LOOP_for_for_for_asn_4153 , CONVOLUTION_LOOP_for_for_for_asn_4155});
  assign COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4145
      , CONVOLUTION_LOOP_for_for_for_asn_4147 , CONVOLUTION_LOOP_for_for_for_asn_4149});
  assign COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4139
      , CONVOLUTION_LOOP_for_for_for_asn_4141 , CONVOLUTION_LOOP_for_for_for_asn_4143});
  assign COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4133
      , CONVOLUTION_LOOP_for_for_for_asn_4135 , CONVOLUTION_LOOP_for_for_for_asn_4137});
  assign COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4127
      , CONVOLUTION_LOOP_for_for_for_asn_4129 , CONVOLUTION_LOOP_for_for_for_asn_4131});
  assign COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4121
      , CONVOLUTION_LOOP_for_for_for_asn_4123 , CONVOLUTION_LOOP_for_for_for_asn_4125});
  assign COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4115
      , CONVOLUTION_LOOP_for_for_for_asn_4117 , CONVOLUTION_LOOP_for_for_for_asn_4119});
  assign COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4109
      , CONVOLUTION_LOOP_for_for_for_asn_4111 , CONVOLUTION_LOOP_for_for_for_asn_4113});
  assign COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4103
      , CONVOLUTION_LOOP_for_for_for_asn_4105 , CONVOLUTION_LOOP_for_for_for_asn_4107});
  assign COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4097
      , CONVOLUTION_LOOP_for_for_for_asn_4099 , CONVOLUTION_LOOP_for_for_for_asn_4101});
  assign COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4091
      , CONVOLUTION_LOOP_for_for_for_asn_4093 , CONVOLUTION_LOOP_for_for_for_asn_4095});
  assign COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4085
      , CONVOLUTION_LOOP_for_for_for_asn_4087 , CONVOLUTION_LOOP_for_for_for_asn_4089});
  assign COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4079
      , CONVOLUTION_LOOP_for_for_for_asn_4081 , CONVOLUTION_LOOP_for_for_for_asn_4083});
  assign COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4073
      , CONVOLUTION_LOOP_for_for_for_asn_4075 , CONVOLUTION_LOOP_for_for_for_asn_4077});
  assign COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4067
      , CONVOLUTION_LOOP_for_for_for_asn_4069 , CONVOLUTION_LOOP_for_for_for_asn_4071});
  assign COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4061
      , CONVOLUTION_LOOP_for_for_for_asn_4063 , CONVOLUTION_LOOP_for_for_for_asn_4065});
  assign COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4055
      , CONVOLUTION_LOOP_for_for_for_asn_4057 , CONVOLUTION_LOOP_for_for_for_asn_4059});
  assign COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4049
      , CONVOLUTION_LOOP_for_for_for_asn_4051 , CONVOLUTION_LOOP_for_for_for_asn_4053});
  assign COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4043
      , CONVOLUTION_LOOP_for_for_for_asn_4045 , CONVOLUTION_LOOP_for_for_for_asn_4047});
  assign COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4037
      , CONVOLUTION_LOOP_for_for_for_asn_4039 , CONVOLUTION_LOOP_for_for_for_asn_4041});
  assign COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4031
      , CONVOLUTION_LOOP_for_for_for_asn_4033 , CONVOLUTION_LOOP_for_for_for_asn_4035});
  assign COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4025
      , CONVOLUTION_LOOP_for_for_for_asn_4027 , CONVOLUTION_LOOP_for_for_for_asn_4029});
  assign COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4019
      , CONVOLUTION_LOOP_for_for_for_asn_4021 , CONVOLUTION_LOOP_for_for_for_asn_4023});
  assign COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4013
      , CONVOLUTION_LOOP_for_for_for_asn_4015 , CONVOLUTION_LOOP_for_for_for_asn_4017});
  assign COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4007
      , CONVOLUTION_LOOP_for_for_for_asn_4009 , CONVOLUTION_LOOP_for_for_for_asn_4011});
  assign COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_4001
      , CONVOLUTION_LOOP_for_for_for_asn_4003 , CONVOLUTION_LOOP_for_for_for_asn_4005});
  assign COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3995
      , CONVOLUTION_LOOP_for_for_for_asn_3997 , CONVOLUTION_LOOP_for_for_for_asn_3999});
  assign COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3989
      , CONVOLUTION_LOOP_for_for_for_asn_3991 , CONVOLUTION_LOOP_for_for_for_asn_3993});
  assign COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3983
      , CONVOLUTION_LOOP_for_for_for_asn_3985 , CONVOLUTION_LOOP_for_for_for_asn_3987});
  assign COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3977
      , CONVOLUTION_LOOP_for_for_for_asn_3979 , CONVOLUTION_LOOP_for_for_for_asn_3981});
  assign COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3971
      , CONVOLUTION_LOOP_for_for_for_asn_3973 , CONVOLUTION_LOOP_for_for_for_asn_3975});
  assign COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3965
      , CONVOLUTION_LOOP_for_for_for_asn_3967 , CONVOLUTION_LOOP_for_for_for_asn_3969});
  assign COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3959
      , CONVOLUTION_LOOP_for_for_for_asn_3961 , CONVOLUTION_LOOP_for_for_for_asn_3963});
  assign COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3953
      , CONVOLUTION_LOOP_for_for_for_asn_3955 , CONVOLUTION_LOOP_for_for_for_asn_3957});
  assign COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3947
      , CONVOLUTION_LOOP_for_for_for_asn_3949 , CONVOLUTION_LOOP_for_for_for_asn_3951});
  assign COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3941
      , CONVOLUTION_LOOP_for_for_for_asn_3943 , CONVOLUTION_LOOP_for_for_for_asn_3945});
  assign COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3935
      , CONVOLUTION_LOOP_for_for_for_asn_3937 , CONVOLUTION_LOOP_for_for_for_asn_3939});
  assign COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3929
      , CONVOLUTION_LOOP_for_for_for_asn_3931 , CONVOLUTION_LOOP_for_for_for_asn_3933});
  assign COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3923
      , CONVOLUTION_LOOP_for_for_for_asn_3925 , CONVOLUTION_LOOP_for_for_for_asn_3927});
  assign COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3917
      , CONVOLUTION_LOOP_for_for_for_asn_3919 , CONVOLUTION_LOOP_for_for_for_asn_3921});
  assign COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3911
      , CONVOLUTION_LOOP_for_for_for_asn_3913 , CONVOLUTION_LOOP_for_for_for_asn_3915});
  assign COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3905
      , CONVOLUTION_LOOP_for_for_for_asn_3907 , CONVOLUTION_LOOP_for_for_for_asn_3909});
  assign COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3899
      , CONVOLUTION_LOOP_for_for_for_asn_3901 , CONVOLUTION_LOOP_for_for_for_asn_3903});
  assign COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3893
      , CONVOLUTION_LOOP_for_for_for_asn_3895 , CONVOLUTION_LOOP_for_for_for_asn_3897});
  assign COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3887
      , CONVOLUTION_LOOP_for_for_for_asn_3889 , CONVOLUTION_LOOP_for_for_for_asn_3891});
  assign COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3881
      , CONVOLUTION_LOOP_for_for_for_asn_3883 , CONVOLUTION_LOOP_for_for_for_asn_3885});
  assign COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3875
      , CONVOLUTION_LOOP_for_for_for_asn_3877 , CONVOLUTION_LOOP_for_for_for_asn_3879});
  assign COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3869
      , CONVOLUTION_LOOP_for_for_for_asn_3871 , CONVOLUTION_LOOP_for_for_for_asn_3873});
  assign COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3863
      , CONVOLUTION_LOOP_for_for_for_asn_3865 , CONVOLUTION_LOOP_for_for_for_asn_3867});
  assign COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3857
      , CONVOLUTION_LOOP_for_for_for_asn_3859 , CONVOLUTION_LOOP_for_for_for_asn_3861});
  assign COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3851
      , CONVOLUTION_LOOP_for_for_for_asn_3853 , CONVOLUTION_LOOP_for_for_for_asn_3855});
  assign COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3845
      , CONVOLUTION_LOOP_for_for_for_asn_3847 , CONVOLUTION_LOOP_for_for_for_asn_3849});
  assign COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3839
      , CONVOLUTION_LOOP_for_for_for_asn_3841 , CONVOLUTION_LOOP_for_for_for_asn_3843});
  assign COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3833
      , CONVOLUTION_LOOP_for_for_for_asn_3835 , CONVOLUTION_LOOP_for_for_for_asn_3837});
  assign COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3827
      , CONVOLUTION_LOOP_for_for_for_asn_3829 , CONVOLUTION_LOOP_for_for_for_asn_3831});
  assign COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3821
      , CONVOLUTION_LOOP_for_for_for_asn_3823 , CONVOLUTION_LOOP_for_for_for_asn_3825});
  assign COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3815
      , CONVOLUTION_LOOP_for_for_for_asn_3817 , CONVOLUTION_LOOP_for_for_for_asn_3819});
  assign COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3809
      , CONVOLUTION_LOOP_for_for_for_asn_3811 , CONVOLUTION_LOOP_for_for_for_asn_3813});
  assign COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3803
      , CONVOLUTION_LOOP_for_for_for_asn_3805 , CONVOLUTION_LOOP_for_for_for_asn_3807});
  assign COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3797
      , CONVOLUTION_LOOP_for_for_for_asn_3799 , CONVOLUTION_LOOP_for_for_for_asn_3801});
  assign COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3791
      , CONVOLUTION_LOOP_for_for_for_asn_3793 , CONVOLUTION_LOOP_for_for_for_asn_3795});
  assign COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3785
      , CONVOLUTION_LOOP_for_for_for_asn_3787 , CONVOLUTION_LOOP_for_for_for_asn_3789});
  assign COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3779
      , CONVOLUTION_LOOP_for_for_for_asn_3781 , CONVOLUTION_LOOP_for_for_for_asn_3783});
  assign COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3773
      , CONVOLUTION_LOOP_for_for_for_asn_3775 , CONVOLUTION_LOOP_for_for_for_asn_3777});
  assign COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3767
      , CONVOLUTION_LOOP_for_for_for_asn_3769 , CONVOLUTION_LOOP_for_for_for_asn_3771});
  assign COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3761
      , CONVOLUTION_LOOP_for_for_for_asn_3763 , CONVOLUTION_LOOP_for_for_for_asn_3765});
  assign COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3755
      , CONVOLUTION_LOOP_for_for_for_asn_3757 , CONVOLUTION_LOOP_for_for_for_asn_3759});
  assign COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3749
      , CONVOLUTION_LOOP_for_for_for_asn_3751 , CONVOLUTION_LOOP_for_for_for_asn_3753});
  assign COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3743
      , CONVOLUTION_LOOP_for_for_for_asn_3745 , CONVOLUTION_LOOP_for_for_for_asn_3747});
  assign COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3737
      , CONVOLUTION_LOOP_for_for_for_asn_3739 , CONVOLUTION_LOOP_for_for_for_asn_3741});
  assign COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3731
      , CONVOLUTION_LOOP_for_for_for_asn_3733 , CONVOLUTION_LOOP_for_for_for_asn_3735});
  assign COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3725
      , CONVOLUTION_LOOP_for_for_for_asn_3727 , CONVOLUTION_LOOP_for_for_for_asn_3729});
  assign COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3719
      , CONVOLUTION_LOOP_for_for_for_asn_3721 , CONVOLUTION_LOOP_for_for_for_asn_3723});
  assign COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3713
      , CONVOLUTION_LOOP_for_for_for_asn_3715 , CONVOLUTION_LOOP_for_for_for_asn_3717});
  assign COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3707
      , CONVOLUTION_LOOP_for_for_for_asn_3709 , CONVOLUTION_LOOP_for_for_for_asn_3711});
  assign COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3701
      , CONVOLUTION_LOOP_for_for_for_asn_3703 , CONVOLUTION_LOOP_for_for_for_asn_3705});
  assign COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3695
      , CONVOLUTION_LOOP_for_for_for_asn_3697 , CONVOLUTION_LOOP_for_for_for_asn_3699});
  assign COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3689
      , CONVOLUTION_LOOP_for_for_for_asn_3691 , CONVOLUTION_LOOP_for_for_for_asn_3693});
  assign COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3683
      , CONVOLUTION_LOOP_for_for_for_asn_3685 , CONVOLUTION_LOOP_for_for_for_asn_3687});
  assign COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3677
      , CONVOLUTION_LOOP_for_for_for_asn_3679 , CONVOLUTION_LOOP_for_for_for_asn_3681});
  assign COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3671
      , CONVOLUTION_LOOP_for_for_for_asn_3673 , CONVOLUTION_LOOP_for_for_for_asn_3675});
  assign COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3665
      , CONVOLUTION_LOOP_for_for_for_asn_3667 , CONVOLUTION_LOOP_for_for_for_asn_3669});
  assign COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3659
      , CONVOLUTION_LOOP_for_for_for_asn_3661 , CONVOLUTION_LOOP_for_for_for_asn_3663});
  assign COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3653
      , CONVOLUTION_LOOP_for_for_for_asn_3655 , CONVOLUTION_LOOP_for_for_for_asn_3657});
  assign COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3647
      , CONVOLUTION_LOOP_for_for_for_asn_3649 , CONVOLUTION_LOOP_for_for_for_asn_3651});
  assign COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3641
      , CONVOLUTION_LOOP_for_for_for_asn_3643 , CONVOLUTION_LOOP_for_for_for_asn_3645});
  assign COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3635
      , CONVOLUTION_LOOP_for_for_for_asn_3637 , CONVOLUTION_LOOP_for_for_for_asn_3639});
  assign COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3629
      , CONVOLUTION_LOOP_for_for_for_asn_3631 , CONVOLUTION_LOOP_for_for_for_asn_3633});
  assign COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3623
      , CONVOLUTION_LOOP_for_for_for_asn_3625 , CONVOLUTION_LOOP_for_for_for_asn_3627});
  assign COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3617
      , CONVOLUTION_LOOP_for_for_for_asn_3619 , CONVOLUTION_LOOP_for_for_for_asn_3621});
  assign COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3611
      , CONVOLUTION_LOOP_for_for_for_asn_3613 , CONVOLUTION_LOOP_for_for_for_asn_3615});
  assign COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3605
      , CONVOLUTION_LOOP_for_for_for_asn_3607 , CONVOLUTION_LOOP_for_for_for_asn_3609});
  assign COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3599
      , CONVOLUTION_LOOP_for_for_for_asn_3601 , CONVOLUTION_LOOP_for_for_for_asn_3603});
  assign COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3593
      , CONVOLUTION_LOOP_for_for_for_asn_3595 , CONVOLUTION_LOOP_for_for_for_asn_3597});
  assign COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3587
      , CONVOLUTION_LOOP_for_for_for_asn_3589 , CONVOLUTION_LOOP_for_for_for_asn_3591});
  assign COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3581
      , CONVOLUTION_LOOP_for_for_for_asn_3583 , CONVOLUTION_LOOP_for_for_for_asn_3585});
  assign COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_3 = MUX1HOT_v_11_3_2(COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_2,
      ({{10{CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}}, CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0}),
      ({CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      , (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[54:45])}), {CONVOLUTION_LOOP_for_for_for_asn_3575
      , CONVOLUTION_LOOP_for_for_for_asn_3577 , CONVOLUTION_LOOP_for_for_for_asn_3579});
  assign COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5513 , CONVOLUTION_LOOP_for_for_for_asn_5515
      , CONVOLUTION_LOOP_for_for_for_asn_5517});
  assign COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5507 , CONVOLUTION_LOOP_for_for_for_asn_5509
      , CONVOLUTION_LOOP_for_for_for_asn_5511});
  assign COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5501 , CONVOLUTION_LOOP_for_for_for_asn_5503
      , CONVOLUTION_LOOP_for_for_for_asn_5505});
  assign COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5495 , CONVOLUTION_LOOP_for_for_for_asn_5497
      , CONVOLUTION_LOOP_for_for_for_asn_5499});
  assign COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5489 , CONVOLUTION_LOOP_for_for_for_asn_5491
      , CONVOLUTION_LOOP_for_for_for_asn_5493});
  assign COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5483 , CONVOLUTION_LOOP_for_for_for_asn_5485
      , CONVOLUTION_LOOP_for_for_for_asn_5487});
  assign COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5477 , CONVOLUTION_LOOP_for_for_for_asn_5479
      , CONVOLUTION_LOOP_for_for_for_asn_5481});
  assign COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5471 , CONVOLUTION_LOOP_for_for_for_asn_5473
      , CONVOLUTION_LOOP_for_for_for_asn_5475});
  assign COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5465 , CONVOLUTION_LOOP_for_for_for_asn_5467
      , CONVOLUTION_LOOP_for_for_for_asn_5469});
  assign COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5459 , CONVOLUTION_LOOP_for_for_for_asn_5461
      , CONVOLUTION_LOOP_for_for_for_asn_5463});
  assign COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5453 , CONVOLUTION_LOOP_for_for_for_asn_5455
      , CONVOLUTION_LOOP_for_for_for_asn_5457});
  assign COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5447 , CONVOLUTION_LOOP_for_for_for_asn_5449
      , CONVOLUTION_LOOP_for_for_for_asn_5451});
  assign COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5441 , CONVOLUTION_LOOP_for_for_for_asn_5443
      , CONVOLUTION_LOOP_for_for_for_asn_5445});
  assign COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5435 , CONVOLUTION_LOOP_for_for_for_asn_5437
      , CONVOLUTION_LOOP_for_for_for_asn_5439});
  assign COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5429 , CONVOLUTION_LOOP_for_for_for_asn_5431
      , CONVOLUTION_LOOP_for_for_for_asn_5433});
  assign COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5423 , CONVOLUTION_LOOP_for_for_for_asn_5425
      , CONVOLUTION_LOOP_for_for_for_asn_5427});
  assign COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5417 , CONVOLUTION_LOOP_for_for_for_asn_5419
      , CONVOLUTION_LOOP_for_for_for_asn_5421});
  assign COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5411 , CONVOLUTION_LOOP_for_for_for_asn_5413
      , CONVOLUTION_LOOP_for_for_for_asn_5415});
  assign COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5405 , CONVOLUTION_LOOP_for_for_for_asn_5407
      , CONVOLUTION_LOOP_for_for_for_asn_5409});
  assign COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5399 , CONVOLUTION_LOOP_for_for_for_asn_5401
      , CONVOLUTION_LOOP_for_for_for_asn_5403});
  assign COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5393 , CONVOLUTION_LOOP_for_for_for_asn_5395
      , CONVOLUTION_LOOP_for_for_for_asn_5397});
  assign COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5387 , CONVOLUTION_LOOP_for_for_for_asn_5389
      , CONVOLUTION_LOOP_for_for_for_asn_5391});
  assign COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5381 , CONVOLUTION_LOOP_for_for_for_asn_5383
      , CONVOLUTION_LOOP_for_for_for_asn_5385});
  assign COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5375 , CONVOLUTION_LOOP_for_for_for_asn_5377
      , CONVOLUTION_LOOP_for_for_for_asn_5379});
  assign COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5369 , CONVOLUTION_LOOP_for_for_for_asn_5371
      , CONVOLUTION_LOOP_for_for_for_asn_5373});
  assign COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5363 , CONVOLUTION_LOOP_for_for_for_asn_5365
      , CONVOLUTION_LOOP_for_for_for_asn_5367});
  assign COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5357 , CONVOLUTION_LOOP_for_for_for_asn_5359
      , CONVOLUTION_LOOP_for_for_for_asn_5361});
  assign COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5351 , CONVOLUTION_LOOP_for_for_for_asn_5353
      , CONVOLUTION_LOOP_for_for_for_asn_5355});
  assign COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5345 , CONVOLUTION_LOOP_for_for_for_asn_5347
      , CONVOLUTION_LOOP_for_for_for_asn_5349});
  assign COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5339 , CONVOLUTION_LOOP_for_for_for_asn_5341
      , CONVOLUTION_LOOP_for_for_for_asn_5343});
  assign COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5333 , CONVOLUTION_LOOP_for_for_for_asn_5335
      , CONVOLUTION_LOOP_for_for_for_asn_5337});
  assign COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5327 , CONVOLUTION_LOOP_for_for_for_asn_5329
      , CONVOLUTION_LOOP_for_for_for_asn_5331});
  assign COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5321 , CONVOLUTION_LOOP_for_for_for_asn_5323
      , CONVOLUTION_LOOP_for_for_for_asn_5325});
  assign COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5315 , CONVOLUTION_LOOP_for_for_for_asn_5317
      , CONVOLUTION_LOOP_for_for_for_asn_5319});
  assign COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5309 , CONVOLUTION_LOOP_for_for_for_asn_5311
      , CONVOLUTION_LOOP_for_for_for_asn_5313});
  assign COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5303 , CONVOLUTION_LOOP_for_for_for_asn_5305
      , CONVOLUTION_LOOP_for_for_for_asn_5307});
  assign COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5297 , CONVOLUTION_LOOP_for_for_for_asn_5299
      , CONVOLUTION_LOOP_for_for_for_asn_5301});
  assign COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5291 , CONVOLUTION_LOOP_for_for_for_asn_5293
      , CONVOLUTION_LOOP_for_for_for_asn_5295});
  assign COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5285 , CONVOLUTION_LOOP_for_for_for_asn_5287
      , CONVOLUTION_LOOP_for_for_for_asn_5289});
  assign COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5279 , CONVOLUTION_LOOP_for_for_for_asn_5281
      , CONVOLUTION_LOOP_for_for_for_asn_5283});
  assign COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5273 , CONVOLUTION_LOOP_for_for_for_asn_5275
      , CONVOLUTION_LOOP_for_for_for_asn_5277});
  assign COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5267 , CONVOLUTION_LOOP_for_for_for_asn_5269
      , CONVOLUTION_LOOP_for_for_for_asn_5271});
  assign COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5261 , CONVOLUTION_LOOP_for_for_for_asn_5263
      , CONVOLUTION_LOOP_for_for_for_asn_5265});
  assign COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5255 , CONVOLUTION_LOOP_for_for_for_asn_5257
      , CONVOLUTION_LOOP_for_for_for_asn_5259});
  assign COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5249 , CONVOLUTION_LOOP_for_for_for_asn_5251
      , CONVOLUTION_LOOP_for_for_for_asn_5253});
  assign COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5243 , CONVOLUTION_LOOP_for_for_for_asn_5245
      , CONVOLUTION_LOOP_for_for_for_asn_5247});
  assign COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5237 , CONVOLUTION_LOOP_for_for_for_asn_5239
      , CONVOLUTION_LOOP_for_for_for_asn_5241});
  assign COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5231 , CONVOLUTION_LOOP_for_for_for_asn_5233
      , CONVOLUTION_LOOP_for_for_for_asn_5235});
  assign COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5225 , CONVOLUTION_LOOP_for_for_for_asn_5227
      , CONVOLUTION_LOOP_for_for_for_asn_5229});
  assign COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5219 , CONVOLUTION_LOOP_for_for_for_asn_5221
      , CONVOLUTION_LOOP_for_for_for_asn_5223});
  assign COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5213 , CONVOLUTION_LOOP_for_for_for_asn_5215
      , CONVOLUTION_LOOP_for_for_for_asn_5217});
  assign COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5207 , CONVOLUTION_LOOP_for_for_for_asn_5209
      , CONVOLUTION_LOOP_for_for_for_asn_5211});
  assign COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5201 , CONVOLUTION_LOOP_for_for_for_asn_5203
      , CONVOLUTION_LOOP_for_for_for_asn_5205});
  assign COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5195 , CONVOLUTION_LOOP_for_for_for_asn_5197
      , CONVOLUTION_LOOP_for_for_for_asn_5199});
  assign COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5189 , CONVOLUTION_LOOP_for_for_for_asn_5191
      , CONVOLUTION_LOOP_for_for_for_asn_5193});
  assign COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5183 , CONVOLUTION_LOOP_for_for_for_asn_5185
      , CONVOLUTION_LOOP_for_for_for_asn_5187});
  assign COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5177 , CONVOLUTION_LOOP_for_for_for_asn_5179
      , CONVOLUTION_LOOP_for_for_for_asn_5181});
  assign COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5171 , CONVOLUTION_LOOP_for_for_for_asn_5173
      , CONVOLUTION_LOOP_for_for_for_asn_5175});
  assign COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5165 , CONVOLUTION_LOOP_for_for_for_asn_5167
      , CONVOLUTION_LOOP_for_for_for_asn_5169});
  assign COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5159 , CONVOLUTION_LOOP_for_for_for_asn_5161
      , CONVOLUTION_LOOP_for_for_for_asn_5163});
  assign COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5153 , CONVOLUTION_LOOP_for_for_for_asn_5155
      , CONVOLUTION_LOOP_for_for_for_asn_5157});
  assign COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5147 , CONVOLUTION_LOOP_for_for_for_asn_5149
      , CONVOLUTION_LOOP_for_for_for_asn_5151});
  assign COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5141 , CONVOLUTION_LOOP_for_for_for_asn_5143
      , CONVOLUTION_LOOP_for_for_for_asn_5145});
  assign COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5135 , CONVOLUTION_LOOP_for_for_for_asn_5137
      , CONVOLUTION_LOOP_for_for_for_asn_5139});
  assign COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5129 , CONVOLUTION_LOOP_for_for_for_asn_5131
      , CONVOLUTION_LOOP_for_for_for_asn_5133});
  assign COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5123 , CONVOLUTION_LOOP_for_for_for_asn_5125
      , CONVOLUTION_LOOP_for_for_for_asn_5127});
  assign COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5117 , CONVOLUTION_LOOP_for_for_for_asn_5119
      , CONVOLUTION_LOOP_for_for_for_asn_5121});
  assign COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5111 , CONVOLUTION_LOOP_for_for_for_asn_5113
      , CONVOLUTION_LOOP_for_for_for_asn_5115});
  assign COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5105 , CONVOLUTION_LOOP_for_for_for_asn_5107
      , CONVOLUTION_LOOP_for_for_for_asn_5109});
  assign COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5099 , CONVOLUTION_LOOP_for_for_for_asn_5101
      , CONVOLUTION_LOOP_for_for_for_asn_5103});
  assign COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5093 , CONVOLUTION_LOOP_for_for_for_asn_5095
      , CONVOLUTION_LOOP_for_for_for_asn_5097});
  assign COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5087 , CONVOLUTION_LOOP_for_for_for_asn_5089
      , CONVOLUTION_LOOP_for_for_for_asn_5091});
  assign COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5081 , CONVOLUTION_LOOP_for_for_for_asn_5083
      , CONVOLUTION_LOOP_for_for_for_asn_5085});
  assign COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5075 , CONVOLUTION_LOOP_for_for_for_asn_5077
      , CONVOLUTION_LOOP_for_for_for_asn_5079});
  assign COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5069 , CONVOLUTION_LOOP_for_for_for_asn_5071
      , CONVOLUTION_LOOP_for_for_for_asn_5073});
  assign COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5063 , CONVOLUTION_LOOP_for_for_for_asn_5065
      , CONVOLUTION_LOOP_for_for_for_asn_5067});
  assign COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5057 , CONVOLUTION_LOOP_for_for_for_asn_5059
      , CONVOLUTION_LOOP_for_for_for_asn_5061});
  assign COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5051 , CONVOLUTION_LOOP_for_for_for_asn_5053
      , CONVOLUTION_LOOP_for_for_for_asn_5055});
  assign COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5045 , CONVOLUTION_LOOP_for_for_for_asn_5047
      , CONVOLUTION_LOOP_for_for_for_asn_5049});
  assign COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5039 , CONVOLUTION_LOOP_for_for_for_asn_5041
      , CONVOLUTION_LOOP_for_for_for_asn_5043});
  assign COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5033 , CONVOLUTION_LOOP_for_for_for_asn_5035
      , CONVOLUTION_LOOP_for_for_for_asn_5037});
  assign COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5027 , CONVOLUTION_LOOP_for_for_for_asn_5029
      , CONVOLUTION_LOOP_for_for_for_asn_5031});
  assign COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5021 , CONVOLUTION_LOOP_for_for_for_asn_5023
      , CONVOLUTION_LOOP_for_for_for_asn_5025});
  assign COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5015 , CONVOLUTION_LOOP_for_for_for_asn_5017
      , CONVOLUTION_LOOP_for_for_for_asn_5019});
  assign COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5009 , CONVOLUTION_LOOP_for_for_for_asn_5011
      , CONVOLUTION_LOOP_for_for_for_asn_5013});
  assign COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_5003 , CONVOLUTION_LOOP_for_for_for_asn_5005
      , CONVOLUTION_LOOP_for_for_for_asn_5007});
  assign COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4997 , CONVOLUTION_LOOP_for_for_for_asn_4999
      , CONVOLUTION_LOOP_for_for_for_asn_5001});
  assign COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4991 , CONVOLUTION_LOOP_for_for_for_asn_4993
      , CONVOLUTION_LOOP_for_for_for_asn_4995});
  assign COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4985 , CONVOLUTION_LOOP_for_for_for_asn_4987
      , CONVOLUTION_LOOP_for_for_for_asn_4989});
  assign COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4979 , CONVOLUTION_LOOP_for_for_for_asn_4981
      , CONVOLUTION_LOOP_for_for_for_asn_4983});
  assign COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4973 , CONVOLUTION_LOOP_for_for_for_asn_4975
      , CONVOLUTION_LOOP_for_for_for_asn_4977});
  assign COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4967 , CONVOLUTION_LOOP_for_for_for_asn_4969
      , CONVOLUTION_LOOP_for_for_for_asn_4971});
  assign COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4961 , CONVOLUTION_LOOP_for_for_for_asn_4963
      , CONVOLUTION_LOOP_for_for_for_asn_4965});
  assign COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4955 , CONVOLUTION_LOOP_for_for_for_asn_4957
      , CONVOLUTION_LOOP_for_for_for_asn_4959});
  assign COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4949 , CONVOLUTION_LOOP_for_for_for_asn_4951
      , CONVOLUTION_LOOP_for_for_for_asn_4953});
  assign COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4943 , CONVOLUTION_LOOP_for_for_for_asn_4945
      , CONVOLUTION_LOOP_for_for_for_asn_4947});
  assign COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4937 , CONVOLUTION_LOOP_for_for_for_asn_4939
      , CONVOLUTION_LOOP_for_for_for_asn_4941});
  assign COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4931 , CONVOLUTION_LOOP_for_for_for_asn_4933
      , CONVOLUTION_LOOP_for_for_for_asn_4935});
  assign COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4925 , CONVOLUTION_LOOP_for_for_for_asn_4927
      , CONVOLUTION_LOOP_for_for_for_asn_4929});
  assign COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4919 , CONVOLUTION_LOOP_for_for_for_asn_4921
      , CONVOLUTION_LOOP_for_for_for_asn_4923});
  assign COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4913 , CONVOLUTION_LOOP_for_for_for_asn_4915
      , CONVOLUTION_LOOP_for_for_for_asn_4917});
  assign COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4907 , CONVOLUTION_LOOP_for_for_for_asn_4909
      , CONVOLUTION_LOOP_for_for_for_asn_4911});
  assign COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4901 , CONVOLUTION_LOOP_for_for_for_asn_4903
      , CONVOLUTION_LOOP_for_for_for_asn_4905});
  assign COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4895 , CONVOLUTION_LOOP_for_for_for_asn_4897
      , CONVOLUTION_LOOP_for_for_for_asn_4899});
  assign COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4889 , CONVOLUTION_LOOP_for_for_for_asn_4891
      , CONVOLUTION_LOOP_for_for_for_asn_4893});
  assign COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4883 , CONVOLUTION_LOOP_for_for_for_asn_4885
      , CONVOLUTION_LOOP_for_for_for_asn_4887});
  assign COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4877 , CONVOLUTION_LOOP_for_for_for_asn_4879
      , CONVOLUTION_LOOP_for_for_for_asn_4881});
  assign COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4871 , CONVOLUTION_LOOP_for_for_for_asn_4873
      , CONVOLUTION_LOOP_for_for_for_asn_4875});
  assign COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4865 , CONVOLUTION_LOOP_for_for_for_asn_4867
      , CONVOLUTION_LOOP_for_for_for_asn_4869});
  assign COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4859 , CONVOLUTION_LOOP_for_for_for_asn_4861
      , CONVOLUTION_LOOP_for_for_for_asn_4863});
  assign COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4853 , CONVOLUTION_LOOP_for_for_for_asn_4855
      , CONVOLUTION_LOOP_for_for_for_asn_4857});
  assign COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4847 , CONVOLUTION_LOOP_for_for_for_asn_4849
      , CONVOLUTION_LOOP_for_for_for_asn_4851});
  assign COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4841 , CONVOLUTION_LOOP_for_for_for_asn_4843
      , CONVOLUTION_LOOP_for_for_for_asn_4845});
  assign COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4835 , CONVOLUTION_LOOP_for_for_for_asn_4837
      , CONVOLUTION_LOOP_for_for_for_asn_4839});
  assign COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4829 , CONVOLUTION_LOOP_for_for_for_asn_4831
      , CONVOLUTION_LOOP_for_for_for_asn_4833});
  assign COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4823 , CONVOLUTION_LOOP_for_for_for_asn_4825
      , CONVOLUTION_LOOP_for_for_for_asn_4827});
  assign COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4817 , CONVOLUTION_LOOP_for_for_for_asn_4819
      , CONVOLUTION_LOOP_for_for_for_asn_4821});
  assign COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4811 , CONVOLUTION_LOOP_for_for_for_asn_4813
      , CONVOLUTION_LOOP_for_for_for_asn_4815});
  assign COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4805 , CONVOLUTION_LOOP_for_for_for_asn_4807
      , CONVOLUTION_LOOP_for_for_for_asn_4809});
  assign COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4799 , CONVOLUTION_LOOP_for_for_for_asn_4801
      , CONVOLUTION_LOOP_for_for_for_asn_4803});
  assign COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4793 , CONVOLUTION_LOOP_for_for_for_asn_4795
      , CONVOLUTION_LOOP_for_for_for_asn_4797});
  assign COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4787 , CONVOLUTION_LOOP_for_for_for_asn_4789
      , CONVOLUTION_LOOP_for_for_for_asn_4791});
  assign COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4781 , CONVOLUTION_LOOP_for_for_for_asn_4783
      , CONVOLUTION_LOOP_for_for_for_asn_4785});
  assign COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4775 , CONVOLUTION_LOOP_for_for_for_asn_4777
      , CONVOLUTION_LOOP_for_for_for_asn_4779});
  assign COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4769 , CONVOLUTION_LOOP_for_for_for_asn_4771
      , CONVOLUTION_LOOP_for_for_for_asn_4773});
  assign COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4763 , CONVOLUTION_LOOP_for_for_for_asn_4765
      , CONVOLUTION_LOOP_for_for_for_asn_4767});
  assign COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4757 , CONVOLUTION_LOOP_for_for_for_asn_4759
      , CONVOLUTION_LOOP_for_for_for_asn_4761});
  assign COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4751 , CONVOLUTION_LOOP_for_for_for_asn_4753
      , CONVOLUTION_LOOP_for_for_for_asn_4755});
  assign COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4745 , CONVOLUTION_LOOP_for_for_for_asn_4747
      , CONVOLUTION_LOOP_for_for_for_asn_4749});
  assign COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4739 , CONVOLUTION_LOOP_for_for_for_asn_4741
      , CONVOLUTION_LOOP_for_for_for_asn_4743});
  assign COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4733 , CONVOLUTION_LOOP_for_for_for_asn_4735
      , CONVOLUTION_LOOP_for_for_for_asn_4737});
  assign COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4727 , CONVOLUTION_LOOP_for_for_for_asn_4729
      , CONVOLUTION_LOOP_for_for_for_asn_4731});
  assign COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4721 , CONVOLUTION_LOOP_for_for_for_asn_4723
      , CONVOLUTION_LOOP_for_for_for_asn_4725});
  assign COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4715 , CONVOLUTION_LOOP_for_for_for_asn_4717
      , CONVOLUTION_LOOP_for_for_for_asn_4719});
  assign COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4709 , CONVOLUTION_LOOP_for_for_for_asn_4711
      , CONVOLUTION_LOOP_for_for_for_asn_4713});
  assign COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4703 , CONVOLUTION_LOOP_for_for_for_asn_4705
      , CONVOLUTION_LOOP_for_for_for_asn_4707});
  assign COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4697 , CONVOLUTION_LOOP_for_for_for_asn_4699
      , CONVOLUTION_LOOP_for_for_for_asn_4701});
  assign COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4691 , CONVOLUTION_LOOP_for_for_for_asn_4693
      , CONVOLUTION_LOOP_for_for_for_asn_4695});
  assign COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4685 , CONVOLUTION_LOOP_for_for_for_asn_4687
      , CONVOLUTION_LOOP_for_for_for_asn_4689});
  assign COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4679 , CONVOLUTION_LOOP_for_for_for_asn_4681
      , CONVOLUTION_LOOP_for_for_for_asn_4683});
  assign COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4673 , CONVOLUTION_LOOP_for_for_for_asn_4675
      , CONVOLUTION_LOOP_for_for_for_asn_4677});
  assign COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4667 , CONVOLUTION_LOOP_for_for_for_asn_4669
      , CONVOLUTION_LOOP_for_for_for_asn_4671});
  assign COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4661 , CONVOLUTION_LOOP_for_for_for_asn_4663
      , CONVOLUTION_LOOP_for_for_for_asn_4665});
  assign COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4655 , CONVOLUTION_LOOP_for_for_for_asn_4657
      , CONVOLUTION_LOOP_for_for_for_asn_4659});
  assign COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4649 , CONVOLUTION_LOOP_for_for_for_asn_4651
      , CONVOLUTION_LOOP_for_for_for_asn_4653});
  assign COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4643 , CONVOLUTION_LOOP_for_for_for_asn_4645
      , CONVOLUTION_LOOP_for_for_for_asn_4647});
  assign COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4637 , CONVOLUTION_LOOP_for_for_for_asn_4639
      , CONVOLUTION_LOOP_for_for_for_asn_4641});
  assign COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4631 , CONVOLUTION_LOOP_for_for_for_asn_4633
      , CONVOLUTION_LOOP_for_for_for_asn_4635});
  assign COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4625 , CONVOLUTION_LOOP_for_for_for_asn_4627
      , CONVOLUTION_LOOP_for_for_for_asn_4629});
  assign COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4619 , CONVOLUTION_LOOP_for_for_for_asn_4621
      , CONVOLUTION_LOOP_for_for_for_asn_4623});
  assign COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4613 , CONVOLUTION_LOOP_for_for_for_asn_4615
      , CONVOLUTION_LOOP_for_for_for_asn_4617});
  assign COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4607 , CONVOLUTION_LOOP_for_for_for_asn_4609
      , CONVOLUTION_LOOP_for_for_for_asn_4611});
  assign COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4601 , CONVOLUTION_LOOP_for_for_for_asn_4603
      , CONVOLUTION_LOOP_for_for_for_asn_4605});
  assign COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4595 , CONVOLUTION_LOOP_for_for_for_asn_4597
      , CONVOLUTION_LOOP_for_for_for_asn_4599});
  assign COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4589 , CONVOLUTION_LOOP_for_for_for_asn_4591
      , CONVOLUTION_LOOP_for_for_for_asn_4593});
  assign COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4583 , CONVOLUTION_LOOP_for_for_for_asn_4585
      , CONVOLUTION_LOOP_for_for_for_asn_4587});
  assign COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4577 , CONVOLUTION_LOOP_for_for_for_asn_4579
      , CONVOLUTION_LOOP_for_for_for_asn_4581});
  assign COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4571 , CONVOLUTION_LOOP_for_for_for_asn_4573
      , CONVOLUTION_LOOP_for_for_for_asn_4575});
  assign COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4565 , CONVOLUTION_LOOP_for_for_for_asn_4567
      , CONVOLUTION_LOOP_for_for_for_asn_4569});
  assign COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4559 , CONVOLUTION_LOOP_for_for_for_asn_4561
      , CONVOLUTION_LOOP_for_for_for_asn_4563});
  assign COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4553 , CONVOLUTION_LOOP_for_for_for_asn_4555
      , CONVOLUTION_LOOP_for_for_for_asn_4557});
  assign COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4547 , CONVOLUTION_LOOP_for_for_for_asn_4549
      , CONVOLUTION_LOOP_for_for_for_asn_4551});
  assign COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4541 , CONVOLUTION_LOOP_for_for_for_asn_4543
      , CONVOLUTION_LOOP_for_for_for_asn_4545});
  assign COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4535 , CONVOLUTION_LOOP_for_for_for_asn_4537
      , CONVOLUTION_LOOP_for_for_for_asn_4539});
  assign COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4529 , CONVOLUTION_LOOP_for_for_for_asn_4531
      , CONVOLUTION_LOOP_for_for_for_asn_4533});
  assign COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4523 , CONVOLUTION_LOOP_for_for_for_asn_4525
      , CONVOLUTION_LOOP_for_for_for_asn_4527});
  assign COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4517 , CONVOLUTION_LOOP_for_for_for_asn_4519
      , CONVOLUTION_LOOP_for_for_for_asn_4521});
  assign COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4511 , CONVOLUTION_LOOP_for_for_for_asn_4513
      , CONVOLUTION_LOOP_for_for_for_asn_4515});
  assign COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4505 , CONVOLUTION_LOOP_for_for_for_asn_4507
      , CONVOLUTION_LOOP_for_for_for_asn_4509});
  assign COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4499 , CONVOLUTION_LOOP_for_for_for_asn_4501
      , CONVOLUTION_LOOP_for_for_for_asn_4503});
  assign COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4493 , CONVOLUTION_LOOP_for_for_for_asn_4495
      , CONVOLUTION_LOOP_for_for_for_asn_4497});
  assign COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4487 , CONVOLUTION_LOOP_for_for_for_asn_4489
      , CONVOLUTION_LOOP_for_for_for_asn_4491});
  assign COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4481 , CONVOLUTION_LOOP_for_for_for_asn_4483
      , CONVOLUTION_LOOP_for_for_for_asn_4485});
  assign COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4475 , CONVOLUTION_LOOP_for_for_for_asn_4477
      , CONVOLUTION_LOOP_for_for_for_asn_4479});
  assign COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4469 , CONVOLUTION_LOOP_for_for_for_asn_4471
      , CONVOLUTION_LOOP_for_for_for_asn_4473});
  assign COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4463 , CONVOLUTION_LOOP_for_for_for_asn_4465
      , CONVOLUTION_LOOP_for_for_for_asn_4467});
  assign COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4457 , CONVOLUTION_LOOP_for_for_for_asn_4459
      , CONVOLUTION_LOOP_for_for_for_asn_4461});
  assign COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4451 , CONVOLUTION_LOOP_for_for_for_asn_4453
      , CONVOLUTION_LOOP_for_for_for_asn_4455});
  assign COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4445 , CONVOLUTION_LOOP_for_for_for_asn_4447
      , CONVOLUTION_LOOP_for_for_for_asn_4449});
  assign COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4439 , CONVOLUTION_LOOP_for_for_for_asn_4441
      , CONVOLUTION_LOOP_for_for_for_asn_4443});
  assign COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4433 , CONVOLUTION_LOOP_for_for_for_asn_4435
      , CONVOLUTION_LOOP_for_for_for_asn_4437});
  assign COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4427 , CONVOLUTION_LOOP_for_for_for_asn_4429
      , CONVOLUTION_LOOP_for_for_for_asn_4431});
  assign COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4421 , CONVOLUTION_LOOP_for_for_for_asn_4423
      , CONVOLUTION_LOOP_for_for_for_asn_4425});
  assign COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4415 , CONVOLUTION_LOOP_for_for_for_asn_4417
      , CONVOLUTION_LOOP_for_for_for_asn_4419});
  assign COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4409 , CONVOLUTION_LOOP_for_for_for_asn_4411
      , CONVOLUTION_LOOP_for_for_for_asn_4413});
  assign COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4403 , CONVOLUTION_LOOP_for_for_for_asn_4405
      , CONVOLUTION_LOOP_for_for_for_asn_4407});
  assign COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4397 , CONVOLUTION_LOOP_for_for_for_asn_4399
      , CONVOLUTION_LOOP_for_for_for_asn_4401});
  assign COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4391 , CONVOLUTION_LOOP_for_for_for_asn_4393
      , CONVOLUTION_LOOP_for_for_for_asn_4395});
  assign COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4385 , CONVOLUTION_LOOP_for_for_for_asn_4387
      , CONVOLUTION_LOOP_for_for_for_asn_4389});
  assign COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4379 , CONVOLUTION_LOOP_for_for_for_asn_4381
      , CONVOLUTION_LOOP_for_for_for_asn_4383});
  assign COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4373 , CONVOLUTION_LOOP_for_for_for_asn_4375
      , CONVOLUTION_LOOP_for_for_for_asn_4377});
  assign COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4367 , CONVOLUTION_LOOP_for_for_for_asn_4369
      , CONVOLUTION_LOOP_for_for_for_asn_4371});
  assign COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4361 , CONVOLUTION_LOOP_for_for_for_asn_4363
      , CONVOLUTION_LOOP_for_for_for_asn_4365});
  assign COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4355 , CONVOLUTION_LOOP_for_for_for_asn_4357
      , CONVOLUTION_LOOP_for_for_for_asn_4359});
  assign COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4349 , CONVOLUTION_LOOP_for_for_for_asn_4351
      , CONVOLUTION_LOOP_for_for_for_asn_4353});
  assign COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4343 , CONVOLUTION_LOOP_for_for_for_asn_4345
      , CONVOLUTION_LOOP_for_for_for_asn_4347});
  assign COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4337 , CONVOLUTION_LOOP_for_for_for_asn_4339
      , CONVOLUTION_LOOP_for_for_for_asn_4341});
  assign COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4331 , CONVOLUTION_LOOP_for_for_for_asn_4333
      , CONVOLUTION_LOOP_for_for_for_asn_4335});
  assign COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4325 , CONVOLUTION_LOOP_for_for_for_asn_4327
      , CONVOLUTION_LOOP_for_for_for_asn_4329});
  assign COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4319 , CONVOLUTION_LOOP_for_for_for_asn_4321
      , CONVOLUTION_LOOP_for_for_for_asn_4323});
  assign COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4313 , CONVOLUTION_LOOP_for_for_for_asn_4315
      , CONVOLUTION_LOOP_for_for_for_asn_4317});
  assign COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4307 , CONVOLUTION_LOOP_for_for_for_asn_4309
      , CONVOLUTION_LOOP_for_for_for_asn_4311});
  assign COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4301 , CONVOLUTION_LOOP_for_for_for_asn_4303
      , CONVOLUTION_LOOP_for_for_for_asn_4305});
  assign COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4295 , CONVOLUTION_LOOP_for_for_for_asn_4297
      , CONVOLUTION_LOOP_for_for_for_asn_4299});
  assign COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4289 , CONVOLUTION_LOOP_for_for_for_asn_4291
      , CONVOLUTION_LOOP_for_for_for_asn_4293});
  assign COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4283 , CONVOLUTION_LOOP_for_for_for_asn_4285
      , CONVOLUTION_LOOP_for_for_for_asn_4287});
  assign COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4277 , CONVOLUTION_LOOP_for_for_for_asn_4279
      , CONVOLUTION_LOOP_for_for_for_asn_4281});
  assign COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4271 , CONVOLUTION_LOOP_for_for_for_asn_4273
      , CONVOLUTION_LOOP_for_for_for_asn_4275});
  assign COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4265 , CONVOLUTION_LOOP_for_for_for_asn_4267
      , CONVOLUTION_LOOP_for_for_for_asn_4269});
  assign COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4259 , CONVOLUTION_LOOP_for_for_for_asn_4261
      , CONVOLUTION_LOOP_for_for_for_asn_4263});
  assign COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4253 , CONVOLUTION_LOOP_for_for_for_asn_4255
      , CONVOLUTION_LOOP_for_for_for_asn_4257});
  assign COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4247 , CONVOLUTION_LOOP_for_for_for_asn_4249
      , CONVOLUTION_LOOP_for_for_for_asn_4251});
  assign COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4241 , CONVOLUTION_LOOP_for_for_for_asn_4243
      , CONVOLUTION_LOOP_for_for_for_asn_4245});
  assign COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4235 , CONVOLUTION_LOOP_for_for_for_asn_4237
      , CONVOLUTION_LOOP_for_for_for_asn_4239});
  assign COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4229 , CONVOLUTION_LOOP_for_for_for_asn_4231
      , CONVOLUTION_LOOP_for_for_for_asn_4233});
  assign COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4223 , CONVOLUTION_LOOP_for_for_for_asn_4225
      , CONVOLUTION_LOOP_for_for_for_asn_4227});
  assign COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4217 , CONVOLUTION_LOOP_for_for_for_asn_4219
      , CONVOLUTION_LOOP_for_for_for_asn_4221});
  assign COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4211 , CONVOLUTION_LOOP_for_for_for_asn_4213
      , CONVOLUTION_LOOP_for_for_for_asn_4215});
  assign COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4205 , CONVOLUTION_LOOP_for_for_for_asn_4207
      , CONVOLUTION_LOOP_for_for_for_asn_4209});
  assign COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4199 , CONVOLUTION_LOOP_for_for_for_asn_4201
      , CONVOLUTION_LOOP_for_for_for_asn_4203});
  assign COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4193 , CONVOLUTION_LOOP_for_for_for_asn_4195
      , CONVOLUTION_LOOP_for_for_for_asn_4197});
  assign COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4187 , CONVOLUTION_LOOP_for_for_for_asn_4189
      , CONVOLUTION_LOOP_for_for_for_asn_4191});
  assign COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4181 , CONVOLUTION_LOOP_for_for_for_asn_4183
      , CONVOLUTION_LOOP_for_for_for_asn_4185});
  assign COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4175 , CONVOLUTION_LOOP_for_for_for_asn_4177
      , CONVOLUTION_LOOP_for_for_for_asn_4179});
  assign COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4169 , CONVOLUTION_LOOP_for_for_for_asn_4171
      , CONVOLUTION_LOOP_for_for_for_asn_4173});
  assign COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4163 , CONVOLUTION_LOOP_for_for_for_asn_4165
      , CONVOLUTION_LOOP_for_for_for_asn_4167});
  assign COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4157 , CONVOLUTION_LOOP_for_for_for_asn_4159
      , CONVOLUTION_LOOP_for_for_for_asn_4161});
  assign COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4151 , CONVOLUTION_LOOP_for_for_for_asn_4153
      , CONVOLUTION_LOOP_for_for_for_asn_4155});
  assign COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4145 , CONVOLUTION_LOOP_for_for_for_asn_4147
      , CONVOLUTION_LOOP_for_for_for_asn_4149});
  assign COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4139 , CONVOLUTION_LOOP_for_for_for_asn_4141
      , CONVOLUTION_LOOP_for_for_for_asn_4143});
  assign COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4133 , CONVOLUTION_LOOP_for_for_for_asn_4135
      , CONVOLUTION_LOOP_for_for_for_asn_4137});
  assign COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4127 , CONVOLUTION_LOOP_for_for_for_asn_4129
      , CONVOLUTION_LOOP_for_for_for_asn_4131});
  assign COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4121 , CONVOLUTION_LOOP_for_for_for_asn_4123
      , CONVOLUTION_LOOP_for_for_for_asn_4125});
  assign COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4115 , CONVOLUTION_LOOP_for_for_for_asn_4117
      , CONVOLUTION_LOOP_for_for_for_asn_4119});
  assign COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4109 , CONVOLUTION_LOOP_for_for_for_asn_4111
      , CONVOLUTION_LOOP_for_for_for_asn_4113});
  assign COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4103 , CONVOLUTION_LOOP_for_for_for_asn_4105
      , CONVOLUTION_LOOP_for_for_for_asn_4107});
  assign COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4097 , CONVOLUTION_LOOP_for_for_for_asn_4099
      , CONVOLUTION_LOOP_for_for_for_asn_4101});
  assign COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4091 , CONVOLUTION_LOOP_for_for_for_asn_4093
      , CONVOLUTION_LOOP_for_for_for_asn_4095});
  assign COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4085 , CONVOLUTION_LOOP_for_for_for_asn_4087
      , CONVOLUTION_LOOP_for_for_for_asn_4089});
  assign COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4079 , CONVOLUTION_LOOP_for_for_for_asn_4081
      , CONVOLUTION_LOOP_for_for_for_asn_4083});
  assign COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4073 , CONVOLUTION_LOOP_for_for_for_asn_4075
      , CONVOLUTION_LOOP_for_for_for_asn_4077});
  assign COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4067 , CONVOLUTION_LOOP_for_for_for_asn_4069
      , CONVOLUTION_LOOP_for_for_for_asn_4071});
  assign COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4061 , CONVOLUTION_LOOP_for_for_for_asn_4063
      , CONVOLUTION_LOOP_for_for_for_asn_4065});
  assign COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4055 , CONVOLUTION_LOOP_for_for_for_asn_4057
      , CONVOLUTION_LOOP_for_for_for_asn_4059});
  assign COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4049 , CONVOLUTION_LOOP_for_for_for_asn_4051
      , CONVOLUTION_LOOP_for_for_for_asn_4053});
  assign COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4043 , CONVOLUTION_LOOP_for_for_for_asn_4045
      , CONVOLUTION_LOOP_for_for_for_asn_4047});
  assign COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4037 , CONVOLUTION_LOOP_for_for_for_asn_4039
      , CONVOLUTION_LOOP_for_for_for_asn_4041});
  assign COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4031 , CONVOLUTION_LOOP_for_for_for_asn_4033
      , CONVOLUTION_LOOP_for_for_for_asn_4035});
  assign COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4025 , CONVOLUTION_LOOP_for_for_for_asn_4027
      , CONVOLUTION_LOOP_for_for_for_asn_4029});
  assign COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4019 , CONVOLUTION_LOOP_for_for_for_asn_4021
      , CONVOLUTION_LOOP_for_for_for_asn_4023});
  assign COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4013 , CONVOLUTION_LOOP_for_for_for_asn_4015
      , CONVOLUTION_LOOP_for_for_for_asn_4017});
  assign COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4007 , CONVOLUTION_LOOP_for_for_for_asn_4009
      , CONVOLUTION_LOOP_for_for_for_asn_4011});
  assign COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_4001 , CONVOLUTION_LOOP_for_for_for_asn_4003
      , CONVOLUTION_LOOP_for_for_for_asn_4005});
  assign COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3995 , CONVOLUTION_LOOP_for_for_for_asn_3997
      , CONVOLUTION_LOOP_for_for_for_asn_3999});
  assign COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3989 , CONVOLUTION_LOOP_for_for_for_asn_3991
      , CONVOLUTION_LOOP_for_for_for_asn_3993});
  assign COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3983 , CONVOLUTION_LOOP_for_for_for_asn_3985
      , CONVOLUTION_LOOP_for_for_for_asn_3987});
  assign COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3977 , CONVOLUTION_LOOP_for_for_for_asn_3979
      , CONVOLUTION_LOOP_for_for_for_asn_3981});
  assign COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3971 , CONVOLUTION_LOOP_for_for_for_asn_3973
      , CONVOLUTION_LOOP_for_for_for_asn_3975});
  assign COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3965 , CONVOLUTION_LOOP_for_for_for_asn_3967
      , CONVOLUTION_LOOP_for_for_for_asn_3969});
  assign COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3959 , CONVOLUTION_LOOP_for_for_for_asn_3961
      , CONVOLUTION_LOOP_for_for_for_asn_3963});
  assign COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3953 , CONVOLUTION_LOOP_for_for_for_asn_3955
      , CONVOLUTION_LOOP_for_for_for_asn_3957});
  assign COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3947 , CONVOLUTION_LOOP_for_for_for_asn_3949
      , CONVOLUTION_LOOP_for_for_for_asn_3951});
  assign COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3941 , CONVOLUTION_LOOP_for_for_for_asn_3943
      , CONVOLUTION_LOOP_for_for_for_asn_3945});
  assign COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3935 , CONVOLUTION_LOOP_for_for_for_asn_3937
      , CONVOLUTION_LOOP_for_for_for_asn_3939});
  assign COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3929 , CONVOLUTION_LOOP_for_for_for_asn_3931
      , CONVOLUTION_LOOP_for_for_for_asn_3933});
  assign COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3923 , CONVOLUTION_LOOP_for_for_for_asn_3925
      , CONVOLUTION_LOOP_for_for_for_asn_3927});
  assign COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3917 , CONVOLUTION_LOOP_for_for_for_asn_3919
      , CONVOLUTION_LOOP_for_for_for_asn_3921});
  assign COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3911 , CONVOLUTION_LOOP_for_for_for_asn_3913
      , CONVOLUTION_LOOP_for_for_for_asn_3915});
  assign COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3905 , CONVOLUTION_LOOP_for_for_for_asn_3907
      , CONVOLUTION_LOOP_for_for_for_asn_3909});
  assign COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3899 , CONVOLUTION_LOOP_for_for_for_asn_3901
      , CONVOLUTION_LOOP_for_for_for_asn_3903});
  assign COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3893 , CONVOLUTION_LOOP_for_for_for_asn_3895
      , CONVOLUTION_LOOP_for_for_for_asn_3897});
  assign COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3887 , CONVOLUTION_LOOP_for_for_for_asn_3889
      , CONVOLUTION_LOOP_for_for_for_asn_3891});
  assign COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3881 , CONVOLUTION_LOOP_for_for_for_asn_3883
      , CONVOLUTION_LOOP_for_for_for_asn_3885});
  assign COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3875 , CONVOLUTION_LOOP_for_for_for_asn_3877
      , CONVOLUTION_LOOP_for_for_for_asn_3879});
  assign COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3869 , CONVOLUTION_LOOP_for_for_for_asn_3871
      , CONVOLUTION_LOOP_for_for_for_asn_3873});
  assign COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3863 , CONVOLUTION_LOOP_for_for_for_asn_3865
      , CONVOLUTION_LOOP_for_for_for_asn_3867});
  assign COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3857 , CONVOLUTION_LOOP_for_for_for_asn_3859
      , CONVOLUTION_LOOP_for_for_for_asn_3861});
  assign COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3851 , CONVOLUTION_LOOP_for_for_for_asn_3853
      , CONVOLUTION_LOOP_for_for_for_asn_3855});
  assign COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3845 , CONVOLUTION_LOOP_for_for_for_asn_3847
      , CONVOLUTION_LOOP_for_for_for_asn_3849});
  assign COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3839 , CONVOLUTION_LOOP_for_for_for_asn_3841
      , CONVOLUTION_LOOP_for_for_for_asn_3843});
  assign COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3833 , CONVOLUTION_LOOP_for_for_for_asn_3835
      , CONVOLUTION_LOOP_for_for_for_asn_3837});
  assign COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3827 , CONVOLUTION_LOOP_for_for_for_asn_3829
      , CONVOLUTION_LOOP_for_for_for_asn_3831});
  assign COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3821 , CONVOLUTION_LOOP_for_for_for_asn_3823
      , CONVOLUTION_LOOP_for_for_for_asn_3825});
  assign COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3815 , CONVOLUTION_LOOP_for_for_for_asn_3817
      , CONVOLUTION_LOOP_for_for_for_asn_3819});
  assign COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3809 , CONVOLUTION_LOOP_for_for_for_asn_3811
      , CONVOLUTION_LOOP_for_for_for_asn_3813});
  assign COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3803 , CONVOLUTION_LOOP_for_for_for_asn_3805
      , CONVOLUTION_LOOP_for_for_for_asn_3807});
  assign COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3797 , CONVOLUTION_LOOP_for_for_for_asn_3799
      , CONVOLUTION_LOOP_for_for_for_asn_3801});
  assign COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3791 , CONVOLUTION_LOOP_for_for_for_asn_3793
      , CONVOLUTION_LOOP_for_for_for_asn_3795});
  assign COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3785 , CONVOLUTION_LOOP_for_for_for_asn_3787
      , CONVOLUTION_LOOP_for_for_for_asn_3789});
  assign COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3779 , CONVOLUTION_LOOP_for_for_for_asn_3781
      , CONVOLUTION_LOOP_for_for_for_asn_3783});
  assign COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3773 , CONVOLUTION_LOOP_for_for_for_asn_3775
      , CONVOLUTION_LOOP_for_for_for_asn_3777});
  assign COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3767 , CONVOLUTION_LOOP_for_for_for_asn_3769
      , CONVOLUTION_LOOP_for_for_for_asn_3771});
  assign COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3761 , CONVOLUTION_LOOP_for_for_for_asn_3763
      , CONVOLUTION_LOOP_for_for_for_asn_3765});
  assign COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3755 , CONVOLUTION_LOOP_for_for_for_asn_3757
      , CONVOLUTION_LOOP_for_for_for_asn_3759});
  assign COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3749 , CONVOLUTION_LOOP_for_for_for_asn_3751
      , CONVOLUTION_LOOP_for_for_for_asn_3753});
  assign COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3743 , CONVOLUTION_LOOP_for_for_for_asn_3745
      , CONVOLUTION_LOOP_for_for_for_asn_3747});
  assign COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3737 , CONVOLUTION_LOOP_for_for_for_asn_3739
      , CONVOLUTION_LOOP_for_for_for_asn_3741});
  assign COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3731 , CONVOLUTION_LOOP_for_for_for_asn_3733
      , CONVOLUTION_LOOP_for_for_for_asn_3735});
  assign COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3725 , CONVOLUTION_LOOP_for_for_for_asn_3727
      , CONVOLUTION_LOOP_for_for_for_asn_3729});
  assign COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3719 , CONVOLUTION_LOOP_for_for_for_asn_3721
      , CONVOLUTION_LOOP_for_for_for_asn_3723});
  assign COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3713 , CONVOLUTION_LOOP_for_for_for_asn_3715
      , CONVOLUTION_LOOP_for_for_for_asn_3717});
  assign COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3707 , CONVOLUTION_LOOP_for_for_for_asn_3709
      , CONVOLUTION_LOOP_for_for_for_asn_3711});
  assign COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3701 , CONVOLUTION_LOOP_for_for_for_asn_3703
      , CONVOLUTION_LOOP_for_for_for_asn_3705});
  assign COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3695 , CONVOLUTION_LOOP_for_for_for_asn_3697
      , CONVOLUTION_LOOP_for_for_for_asn_3699});
  assign COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3689 , CONVOLUTION_LOOP_for_for_for_asn_3691
      , CONVOLUTION_LOOP_for_for_for_asn_3693});
  assign COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3683 , CONVOLUTION_LOOP_for_for_for_asn_3685
      , CONVOLUTION_LOOP_for_for_for_asn_3687});
  assign COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3677 , CONVOLUTION_LOOP_for_for_for_asn_3679
      , CONVOLUTION_LOOP_for_for_for_asn_3681});
  assign COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3671 , CONVOLUTION_LOOP_for_for_for_asn_3673
      , CONVOLUTION_LOOP_for_for_for_asn_3675});
  assign COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3665 , CONVOLUTION_LOOP_for_for_for_asn_3667
      , CONVOLUTION_LOOP_for_for_for_asn_3669});
  assign COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3659 , CONVOLUTION_LOOP_for_for_for_asn_3661
      , CONVOLUTION_LOOP_for_for_for_asn_3663});
  assign COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3653 , CONVOLUTION_LOOP_for_for_for_asn_3655
      , CONVOLUTION_LOOP_for_for_for_asn_3657});
  assign COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3647 , CONVOLUTION_LOOP_for_for_for_asn_3649
      , CONVOLUTION_LOOP_for_for_for_asn_3651});
  assign COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3641 , CONVOLUTION_LOOP_for_for_for_asn_3643
      , CONVOLUTION_LOOP_for_for_for_asn_3645});
  assign COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3635 , CONVOLUTION_LOOP_for_for_for_asn_3637
      , CONVOLUTION_LOOP_for_for_for_asn_3639});
  assign COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3629 , CONVOLUTION_LOOP_for_for_for_asn_3631
      , CONVOLUTION_LOOP_for_for_for_asn_3633});
  assign COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3623 , CONVOLUTION_LOOP_for_for_for_asn_3625
      , CONVOLUTION_LOOP_for_for_for_asn_3627});
  assign COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3617 , CONVOLUTION_LOOP_for_for_for_asn_3619
      , CONVOLUTION_LOOP_for_for_for_asn_3621});
  assign COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3611 , CONVOLUTION_LOOP_for_for_for_asn_3613
      , CONVOLUTION_LOOP_for_for_for_asn_3615});
  assign COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3605 , CONVOLUTION_LOOP_for_for_for_asn_3607
      , CONVOLUTION_LOOP_for_for_for_asn_3609});
  assign COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3599 , CONVOLUTION_LOOP_for_for_for_asn_3601
      , CONVOLUTION_LOOP_for_for_for_asn_3603});
  assign COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3593 , CONVOLUTION_LOOP_for_for_for_asn_3595
      , CONVOLUTION_LOOP_for_for_for_asn_3597});
  assign COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3587 , CONVOLUTION_LOOP_for_for_for_asn_3589
      , CONVOLUTION_LOOP_for_for_for_asn_3591});
  assign COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3581 , CONVOLUTION_LOOP_for_for_for_asn_3583
      , CONVOLUTION_LOOP_for_for_for_asn_3585});
  assign COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_3 = MUX1HOT_v_45_3_2(COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_2,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, (CONVOLUTION_LOOP_for_for_for_else_conc_ctmp_56_1_sva_1_54_0[44:0]),
      {CONVOLUTION_LOOP_for_for_for_asn_3575 , CONVOLUTION_LOOP_for_for_for_asn_3577
      , CONVOLUTION_LOOP_for_for_for_asn_3579});
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_7_nl = (CONVOLUTION_LOOP_for_for_for_for_for_mul_9_sdt_sva_1[15])
      & ((CONVOLUTION_LOOP_for_for_for_for_for_mul_9_sdt_sva_1[14:0]!=15'b000000000000000)
      | (CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1[0]));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1 = CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1
      + conv_u2s_1_49(CONVOLUTION_LOOP_for_for_for_for_for_and_7_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[48:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_and_unfl_sva_1 = (CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[48])
      & (~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[47:46]==2'b11)));
  assign CONVOLUTION_LOOP_for_for_for_for_for_nor_ovfl_sva_1 = ~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[48])
      | (~((CONVOLUTION_LOOP_for_for_for_for_for_acc_6_psp_sva_1[47:46]!=2'b00))));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1 = conv_s2u_47_49({CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
      , CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
      , CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1})
      + conv_s2u_48_49(CONVOLUTION_LOOP_for_for_for_for_for_mul_9_sdt_sva_1[63:16]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_9_psp_sva_1[48:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_9_sdt_sva_1 = conv_s2u_64_64($signed((plm_filters_rsci_q_d_mxwt))
      * $signed((plm_inputs_rsci_q_d_mxwt)));
  assign unequal_tmp_1 = ~((conf_info_rsci_idat_mxwt[7:0]==8'b00000001));
  assign nl_if_acc_4_cse_1 = ({(pad_sva_1[6:0]) , 1'b0}) - (conf_info_rsci_idat_mxwt[31:24]);
  assign if_acc_4_cse_1 = nl_if_acc_4_cse_1[7:0];
  assign operator_43_true_and_nl = (pad_acc_psp_sva_1[16]) & (pad_acc_psp_sva_1[0]);
  assign nl_operator_43_true_operator_43_true_acc_nl = (pad_acc_psp_sva_1[8:1]) +
      conv_u2s_1_8(operator_43_true_and_nl);
  assign operator_43_true_operator_43_true_acc_nl = nl_operator_43_true_operator_43_true_acc_nl[7:0];
  assign nl_pad_sva_1 = $signed(operator_43_true_operator_43_true_acc_nl) * $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[15:8]));
  assign pad_sva_1 = nl_pad_sva_1[7:0];
  assign nl_else_acc_2_psp_sva_1 = conv_u2s_10_11(else_acc_4_cse_1) + conv_s2s_9_11({1'b1
      , (conf_info_rsci_idat_mxwt[47:40])});
  assign else_acc_2_psp_sva_1 = nl_else_acc_2_psp_sva_1[10:0];
  assign nl_else_acc_4_cse_1 = conv_u2u_9_10({pad_sva_1 , 1'b0}) + conv_u2u_8_10(~
      (conf_info_rsci_idat_mxwt[31:24])) + 10'b0000000001;
  assign else_acc_4_cse_1 = nl_else_acc_4_cse_1[9:0];
  assign nl_else_acc_psp_sva_1 = conv_u2s_10_11(else_acc_4_cse_1) + conv_s2s_9_11({1'b1
      , (conf_info_rsci_idat_mxwt[55:48])});
  assign else_acc_psp_sva_1 = nl_else_acc_psp_sva_1[10:0];
  assign nl_pad_acc_2_nl = ({1'b1 , (~ (conf_info_rsci_idat_mxwt[55:48]))}) + conv_u2s_8_9(conf_info_rsci_idat_mxwt[31:24])
      + 9'b000000001;
  assign pad_acc_2_nl = nl_pad_acc_2_nl[8:0];
  assign nl_operator_8_false_acc_nl = conv_u2s_8_9(conf_info_rsci_idat_mxwt[55:48])
      + 9'b111111111;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[8:0];
  assign nl_pad_mul_nl = $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[7:0])) * $signed(operator_8_false_acc_nl);
  assign pad_mul_nl = nl_pad_mul_nl[16:0];
  assign nl_pad_acc_psp_sva_1 = conv_s2s_9_17(pad_acc_2_nl) + pad_mul_nl;
  assign pad_acc_psp_sva_1 = nl_pad_acc_psp_sva_1[16:0];
  assign nl_COMPUTE_LOOP_acc_tmp = conv_u2u_4_5(COMPUTE_LOOP_b_4_0_lpi_1_dfm_3_0_1)
      + 5'b00001;
  assign COMPUTE_LOOP_acc_tmp = nl_COMPUTE_LOOP_acc_tmp[4:0];
  assign COMPUTE_LOOP_not_35_nl = ~ exitL_exit_COMPUTE_LOOP_sva;
  assign COMPUTE_LOOP_b_4_0_lpi_1_dfm_3_0_1 = MUX_v_4_2_2(4'b0000, COMPUTE_LOOP_b_4_0_lpi_1_3_0,
      COMPUTE_LOOP_not_35_nl);
  assign nl_operator_8_false_8_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_231_224_mx0)
      + 9'b111111111;
  assign operator_8_false_8_acc_tmp = nl_operator_8_false_8_acc_tmp[8:0];
  assign nl_CONVOLUTION_LOOP_acc_tmp = conv_u2u_5_6(CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_4_0_1)
      + 6'b000001;
  assign CONVOLUTION_LOOP_acc_tmp = nl_CONVOLUTION_LOOP_acc_tmp[5:0];
  assign CONVOLUTION_LOOP_not_13_nl = ~ COMPUTE_LOOP_COMPUTE_LOOP_or_tmp;
  assign CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_4_0_1 = MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_2_4_0,
      CONVOLUTION_LOOP_not_13_nl);
  assign nl_operator_8_false_7_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_71_64_mx0)
      + 9'b111111111;
  assign operator_8_false_7_acc_tmp = nl_operator_8_false_7_acc_tmp[8:0];
  assign nl_CONVOLUTION_LOOP_for_acc_tmp = conv_u2u_5_6(CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0)
      + 6'b000001;
  assign CONVOLUTION_LOOP_for_acc_tmp = nl_CONVOLUTION_LOOP_for_acc_tmp[5:0];
  assign nl_operator_8_false_3_acc_nl = conv_u2s_4_5(CONVOLUTION_LOOP_for_for_i_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_3_acc_nl = nl_operator_8_false_3_acc_nl[4:0];
  assign operator_8_false_3_acc_itm_4_1 = readslicef_5_1_4(operator_8_false_3_acc_nl);
  assign nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2 = CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6
      + 5'b00001;
  assign CONVOLUTION_LOOP_for_for_i_4_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_i_4_0_sva_2[4:0];
  assign CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6 = MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_4,
      lfst_exit_CONVOLUTION_LOOP_for_1_lpi_1_dfm_1);
  assign nl_operator_8_false_5_acc_tmp = conv_u2s_8_9(n_w_out_lpi_1_dfm_3) + 9'b111111111;
  assign operator_8_false_5_acc_tmp = nl_operator_8_false_5_acc_tmp[8:0];
  assign nl_operator_8_false_4_acc_nl = conv_u2s_4_5(CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2[4:1])
      + 5'b10111;
  assign operator_8_false_4_acc_nl = nl_operator_8_false_4_acc_nl[4:0];
  assign operator_8_false_4_acc_itm_4 = readslicef_5_1_4(operator_8_false_4_acc_nl);
  assign nl_operator_8_false_3_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_135_128_mx0)
      + 9'b111111111;
  assign operator_8_false_3_acc_tmp = nl_operator_8_false_3_acc_tmp[8:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6
      + 5'b00001;
  assign CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2[4:0];
  assign CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6 = MUX_v_5_2_2(5'b00000, CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_4,
      lfst_exit_CONVOLUTION_LOOP_for_for_1_lpi_1_dfm_1);
  assign nl_operator_8_false_4_acc_tmp = conv_u2s_8_9(n_h_out_lpi_1_dfm_3) + 9'b111111111;
  assign operator_8_false_4_acc_tmp = nl_operator_8_false_4_acc_tmp[8:0];
  assign nl_operator_8_false_5_acc_nl = ({1'b1 , CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2})
      + 4'b0001;
  assign operator_8_false_5_acc_nl = nl_operator_8_false_5_acc_nl[3:0];
  assign operator_8_false_5_acc_itm_3_1 = readslicef_4_1_3(operator_8_false_5_acc_nl);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2 = CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_4
      + 3'b001;
  assign CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2[2:0];
  assign CONVOLUTION_LOOP_for_for_for_for_not_24_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_4 = MUX_v_3_2_2(3'b000,
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_2, CONVOLUTION_LOOP_for_for_for_for_not_24_nl);
  assign nl_operator_8_false_1_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_103_96_mx0)
      + 9'b111111111;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[8:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp = ~((operator_8_false_1_acc_tmp[7:3]!=5'b00000));
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2 = CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_5
      + 3'b001;
  assign CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2 = nl_CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2[2:0];
  assign CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_4_nl
      = lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0 & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0);
  assign CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_5 = MUX_v_3_2_2(3'b000,
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_3, CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_4_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp = CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_5
      == (operator_8_false_1_acc_tmp[2:0]);
  assign lfst_exit_CONVOLUTION_LOOP_for_for_1_lpi_1_dfm_1 = (~ exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3)
      & lfst_exit_CONVOLUTION_LOOP_for_1_lpi_1_dfm_1;
  assign lfst_exit_CONVOLUTION_LOOP_for_1_lpi_1_dfm_1 = ~(exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3
      | COMPUTE_LOOP_COMPUTE_LOOP_or_tmp);
  assign and_9_tmp = (conf_info_rsci_bawt | (~ COMPUTE_LOOP_asn_itm)) & or_12_cse_1
      & or_13_cse_1 & or_4_cse_1 & or_5_cse_1 & or_6_cse_1 & or_7_cse_1 & or_8_cse_1
      & or_1_cse_1 & or_2_cse_1 & or_cse_1;
  assign or_12_cse_1 = plm_inputs_rsc_req_obj_bawt | nand_26_cse_1;
  assign or_13_cse_1 = plm_filters_rsc_req_obj_bawt | nand_26_cse_1;
  assign or_4_cse_1 = plm_outputs_rsc_req_obj_bawt | (~(exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_2
      & main_stage_v_2));
  assign or_5_cse_1 = plm_filters_rsci_bawt | (~ main_stage_v_2);
  assign or_6_cse_1 = plm_inputs_rsci_bawt | (~ main_stage_v_2);
  assign or_7_cse_1 = plm_filters_rsc_rls_obj_bawt | nand_15_cse_1;
  assign or_8_cse_1 = plm_inputs_rsc_rls_obj_bawt | nand_15_cse_1;
  assign or_1_cse_1 = plm_outputs_rsci_bawt | (~(CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
      & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_3 & main_stage_v_3));
  assign or_2_cse_1 = plm_outputs_rsc_rls_obj_bawt | (~(exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_3
      & main_stage_v_3));
  assign or_cse_1 = done_rsci_bawt | (~(exit_COMPUTE_LOOP_lpi_1_dfm_2_st_4 & main_stage_v_4));
  assign nand_26_cse_1 = ~(exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_1 & main_stage_v_1);
  assign nand_15_cse_1 = ~(exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_2 & main_stage_v_2);
  assign CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_mx0 = MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1,
      CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_1, and_dcpl_84);
  assign nl_CONVOLUTION_LOOP_for_for_for_x_mul_nl = CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6
      * conf_info_crt_lpi_1_dfm_7_0_mx0;
  assign CONVOLUTION_LOOP_for_for_for_x_mul_nl = nl_CONVOLUTION_LOOP_for_for_for_x_mul_nl[7:0];
  assign CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0 = MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_x_mul_nl,
      CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_1, and_dcpl_84);
  assign nl_CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1 = CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6
      * conf_info_crt_lpi_1_dfm_7_0_mx0;
  assign CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1 = nl_CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1[7:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1 = CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6
      + conv_u2u_4_5(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6[4:1]);
  assign CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1 = nl_CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[4:0];
  assign CONVOLUTION_LOOP_for_for_for_asn_3575 = (~(CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3577 = CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3579 = CONVOLUTION_LOOP_for_for_for_else_and_835_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3581 = (~(CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3583 = CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3585 = CONVOLUTION_LOOP_for_for_for_else_and_833_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3587 = (~(CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3589 = CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3591 = CONVOLUTION_LOOP_for_for_for_else_and_831_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3593 = (~(CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3595 = CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3597 = CONVOLUTION_LOOP_for_for_for_else_and_829_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3599 = (~(CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3601 = CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3603 = CONVOLUTION_LOOP_for_for_for_else_and_827_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3605 = (~(CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3607 = CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3609 = CONVOLUTION_LOOP_for_for_for_else_and_825_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3611 = (~(CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3613 = CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3615 = CONVOLUTION_LOOP_for_for_for_else_and_823_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3617 = (~(CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3619 = CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3621 = CONVOLUTION_LOOP_for_for_for_else_and_821_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3623 = (~(CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3625 = CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3627 = CONVOLUTION_LOOP_for_for_for_else_and_819_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3629 = (~(CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3631 = CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3633 = CONVOLUTION_LOOP_for_for_for_else_and_817_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3635 = (~(CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3637 = CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3639 = CONVOLUTION_LOOP_for_for_for_else_and_815_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3641 = (~(CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3643 = CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3645 = CONVOLUTION_LOOP_for_for_for_else_and_813_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3647 = (~(CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3649 = CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3651 = CONVOLUTION_LOOP_for_for_for_else_and_811_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3653 = (~(CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3655 = CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3657 = CONVOLUTION_LOOP_for_for_for_else_and_809_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3659 = (~(CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3661 = CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3663 = CONVOLUTION_LOOP_for_for_for_else_and_807_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3665 = (~(CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3667 = CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3669 = CONVOLUTION_LOOP_for_for_for_else_and_805_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3671 = (~(CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3673 = CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3675 = CONVOLUTION_LOOP_for_for_for_else_and_803_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3677 = (~(CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3679 = CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3681 = CONVOLUTION_LOOP_for_for_for_else_and_801_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3683 = (~(CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3685 = CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3687 = CONVOLUTION_LOOP_for_for_for_else_and_799_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3689 = (~(CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3691 = CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3693 = CONVOLUTION_LOOP_for_for_for_else_and_797_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3695 = (~(CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3697 = CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3699 = CONVOLUTION_LOOP_for_for_for_else_and_795_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3701 = (~(CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3703 = CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3705 = CONVOLUTION_LOOP_for_for_for_else_and_793_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3707 = (~(CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3709 = CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3711 = CONVOLUTION_LOOP_for_for_for_else_and_791_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3713 = (~(CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3715 = CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3717 = CONVOLUTION_LOOP_for_for_for_else_and_789_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3719 = (~(CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3721 = CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3723 = CONVOLUTION_LOOP_for_for_for_else_and_787_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3725 = (~(CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3727 = CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3729 = CONVOLUTION_LOOP_for_for_for_else_and_785_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3731 = (~(CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3733 = CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3735 = CONVOLUTION_LOOP_for_for_for_else_and_783_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3737 = (~(CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3739 = CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3741 = CONVOLUTION_LOOP_for_for_for_else_and_781_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3743 = (~(CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3745 = CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3747 = CONVOLUTION_LOOP_for_for_for_else_and_779_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3749 = (~(CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3751 = CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3753 = CONVOLUTION_LOOP_for_for_for_else_and_777_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3755 = (~(CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3757 = CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3759 = CONVOLUTION_LOOP_for_for_for_else_and_775_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3761 = (~(CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3763 = CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3765 = CONVOLUTION_LOOP_for_for_for_else_and_773_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3767 = (~(CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3769 = CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3771 = CONVOLUTION_LOOP_for_for_for_else_and_771_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3773 = (~(CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3775 = CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3777 = CONVOLUTION_LOOP_for_for_for_else_and_769_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3779 = (~(CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3781 = CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3783 = CONVOLUTION_LOOP_for_for_for_else_and_767_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3785 = (~(CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3787 = CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3789 = CONVOLUTION_LOOP_for_for_for_else_and_765_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3791 = (~(CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3793 = CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3795 = CONVOLUTION_LOOP_for_for_for_else_and_763_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3797 = (~(CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3799 = CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3801 = CONVOLUTION_LOOP_for_for_for_else_and_761_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3803 = (~(CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3805 = CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3807 = CONVOLUTION_LOOP_for_for_for_else_and_759_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3809 = (~(CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3811 = CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3813 = CONVOLUTION_LOOP_for_for_for_else_and_757_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3815 = (~(CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3817 = CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3819 = CONVOLUTION_LOOP_for_for_for_else_and_755_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3821 = (~(CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3823 = CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3825 = CONVOLUTION_LOOP_for_for_for_else_and_753_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3827 = (~(CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3829 = CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3831 = CONVOLUTION_LOOP_for_for_for_else_and_751_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3833 = (~(CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3835 = CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3837 = CONVOLUTION_LOOP_for_for_for_else_and_749_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3839 = (~(CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3841 = CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3843 = CONVOLUTION_LOOP_for_for_for_else_and_747_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3845 = (~(CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3847 = CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3849 = CONVOLUTION_LOOP_for_for_for_else_and_745_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3851 = (~(CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3853 = CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3855 = CONVOLUTION_LOOP_for_for_for_else_and_743_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3857 = (~(CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3859 = CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3861 = CONVOLUTION_LOOP_for_for_for_else_and_741_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3863 = (~(CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3865 = CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3867 = CONVOLUTION_LOOP_for_for_for_else_and_739_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3869 = (~(CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3871 = CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3873 = CONVOLUTION_LOOP_for_for_for_else_and_737_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3875 = (~(CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3877 = CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3879 = CONVOLUTION_LOOP_for_for_for_else_and_735_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3881 = (~(CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3883 = CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3885 = CONVOLUTION_LOOP_for_for_for_else_and_733_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3887 = (~(CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3889 = CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3891 = CONVOLUTION_LOOP_for_for_for_else_and_731_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3893 = (~(CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3895 = CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3897 = CONVOLUTION_LOOP_for_for_for_else_and_729_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3899 = (~(CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3901 = CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3903 = CONVOLUTION_LOOP_for_for_for_else_and_727_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3905 = (~(CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3907 = CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3909 = CONVOLUTION_LOOP_for_for_for_else_and_725_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3911 = (~(CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3913 = CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3915 = CONVOLUTION_LOOP_for_for_for_else_and_723_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3917 = (~(CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3919 = CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3921 = CONVOLUTION_LOOP_for_for_for_else_and_721_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3923 = (~(CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3925 = CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3927 = CONVOLUTION_LOOP_for_for_for_else_and_719_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3929 = (~(CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3931 = CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3933 = CONVOLUTION_LOOP_for_for_for_else_and_717_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3935 = (~(CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3937 = CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3939 = CONVOLUTION_LOOP_for_for_for_else_and_715_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3941 = (~(CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3943 = CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3945 = CONVOLUTION_LOOP_for_for_for_else_and_713_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3947 = (~(CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3949 = CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3951 = CONVOLUTION_LOOP_for_for_for_else_and_711_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3953 = (~(CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3955 = CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3957 = CONVOLUTION_LOOP_for_for_for_else_and_709_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3959 = (~(CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3961 = CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3963 = CONVOLUTION_LOOP_for_for_for_else_and_707_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3965 = (~(CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3967 = CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3969 = CONVOLUTION_LOOP_for_for_for_else_and_705_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3971 = (~(CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3973 = CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3975 = CONVOLUTION_LOOP_for_for_for_else_and_703_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3977 = (~(CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3979 = CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3981 = CONVOLUTION_LOOP_for_for_for_else_and_701_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3983 = (~(CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3985 = CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3987 = CONVOLUTION_LOOP_for_for_for_else_and_699_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3989 = (~(CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3991 = CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3993 = CONVOLUTION_LOOP_for_for_for_else_and_697_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_3995 = (~(CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3997 = CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_3999 = CONVOLUTION_LOOP_for_for_for_else_and_695_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4001 = (~(CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4003 = CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4005 = CONVOLUTION_LOOP_for_for_for_else_and_693_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4007 = (~(CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4009 = CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4011 = CONVOLUTION_LOOP_for_for_for_else_and_691_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4013 = (~(CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4015 = CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4017 = CONVOLUTION_LOOP_for_for_for_else_and_689_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4019 = (~(CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4021 = CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4023 = CONVOLUTION_LOOP_for_for_for_else_and_687_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4025 = (~(CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4027 = CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4029 = CONVOLUTION_LOOP_for_for_for_else_and_685_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4031 = (~(CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4033 = CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4035 = CONVOLUTION_LOOP_for_for_for_else_and_683_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4037 = (~(CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4039 = CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4041 = CONVOLUTION_LOOP_for_for_for_else_and_681_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4043 = (~(CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4045 = CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4047 = CONVOLUTION_LOOP_for_for_for_else_and_679_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4049 = (~(CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4051 = CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4053 = CONVOLUTION_LOOP_for_for_for_else_and_677_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4055 = (~(CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4057 = CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4059 = CONVOLUTION_LOOP_for_for_for_else_and_675_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4061 = (~(CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4063 = CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4065 = CONVOLUTION_LOOP_for_for_for_else_and_673_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4067 = (~(CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4069 = CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4071 = CONVOLUTION_LOOP_for_for_for_else_and_671_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4073 = (~(CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4075 = CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4077 = CONVOLUTION_LOOP_for_for_for_else_and_669_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4079 = (~(CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4081 = CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4083 = CONVOLUTION_LOOP_for_for_for_else_and_667_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4085 = (~(CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4087 = CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4089 = CONVOLUTION_LOOP_for_for_for_else_and_665_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4091 = (~(CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4093 = CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4095 = CONVOLUTION_LOOP_for_for_for_else_and_663_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4097 = (~(CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4099 = CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4101 = CONVOLUTION_LOOP_for_for_for_else_and_661_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4103 = (~(CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4105 = CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4107 = CONVOLUTION_LOOP_for_for_for_else_and_659_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4109 = (~(CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4111 = CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4113 = CONVOLUTION_LOOP_for_for_for_else_and_657_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4115 = (~(CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4117 = CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4119 = CONVOLUTION_LOOP_for_for_for_else_and_655_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4121 = (~(CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4123 = CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4125 = CONVOLUTION_LOOP_for_for_for_else_and_653_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4127 = (~(CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4129 = CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4131 = CONVOLUTION_LOOP_for_for_for_else_and_651_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4133 = (~(CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4135 = CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4137 = CONVOLUTION_LOOP_for_for_for_else_and_649_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4139 = (~(CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4141 = CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4143 = CONVOLUTION_LOOP_for_for_for_else_and_647_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4145 = (~(CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4147 = CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4149 = CONVOLUTION_LOOP_for_for_for_else_and_645_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4151 = (~(CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4153 = CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4155 = CONVOLUTION_LOOP_for_for_for_else_and_643_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4157 = (~(CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4159 = CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4161 = CONVOLUTION_LOOP_for_for_for_else_and_641_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4163 = (~(CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4165 = CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4167 = CONVOLUTION_LOOP_for_for_for_else_and_639_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4169 = (~(CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4171 = CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4173 = CONVOLUTION_LOOP_for_for_for_else_and_637_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4175 = (~(CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4177 = CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4179 = CONVOLUTION_LOOP_for_for_for_else_and_635_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4181 = (~(CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4183 = CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4185 = CONVOLUTION_LOOP_for_for_for_else_and_633_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4187 = (~(CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4189 = CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4191 = CONVOLUTION_LOOP_for_for_for_else_and_631_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4193 = (~(CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4195 = CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4197 = CONVOLUTION_LOOP_for_for_for_else_and_629_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4199 = (~(CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4201 = CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4203 = CONVOLUTION_LOOP_for_for_for_else_and_627_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4205 = (~(CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4207 = CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4209 = CONVOLUTION_LOOP_for_for_for_else_and_625_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4211 = (~(CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4213 = CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4215 = CONVOLUTION_LOOP_for_for_for_else_and_623_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4217 = (~(CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4219 = CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4221 = CONVOLUTION_LOOP_for_for_for_else_and_621_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4223 = (~(CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4225 = CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4227 = CONVOLUTION_LOOP_for_for_for_else_and_619_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4229 = (~(CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4231 = CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4233 = CONVOLUTION_LOOP_for_for_for_else_and_617_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4235 = (~(CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4237 = CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4239 = CONVOLUTION_LOOP_for_for_for_else_and_615_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4241 = (~(CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4243 = CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4245 = CONVOLUTION_LOOP_for_for_for_else_and_613_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4247 = (~(CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4249 = CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4251 = CONVOLUTION_LOOP_for_for_for_else_and_611_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4253 = (~(CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4255 = CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4257 = CONVOLUTION_LOOP_for_for_for_else_and_609_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4259 = (~(CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4261 = CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4263 = CONVOLUTION_LOOP_for_for_for_else_and_607_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4265 = (~(CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4267 = CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4269 = CONVOLUTION_LOOP_for_for_for_else_and_605_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4271 = (~(CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4273 = CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4275 = CONVOLUTION_LOOP_for_for_for_else_and_603_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4277 = (~(CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4279 = CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4281 = CONVOLUTION_LOOP_for_for_for_else_and_601_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4283 = (~(CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4285 = CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4287 = CONVOLUTION_LOOP_for_for_for_else_and_599_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4289 = (~(CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4291 = CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4293 = CONVOLUTION_LOOP_for_for_for_else_and_597_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4295 = (~(CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4297 = CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4299 = CONVOLUTION_LOOP_for_for_for_else_and_595_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4301 = (~(CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4303 = CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4305 = CONVOLUTION_LOOP_for_for_for_else_and_593_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4307 = (~(CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4309 = CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4311 = CONVOLUTION_LOOP_for_for_for_else_and_591_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4313 = (~(CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4315 = CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4317 = CONVOLUTION_LOOP_for_for_for_else_and_589_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4319 = (~(CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4321 = CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4323 = CONVOLUTION_LOOP_for_for_for_else_and_587_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4325 = (~(CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4327 = CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4329 = CONVOLUTION_LOOP_for_for_for_else_and_585_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4331 = (~(CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4333 = CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4335 = CONVOLUTION_LOOP_for_for_for_else_and_583_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4337 = (~(CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4339 = CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4341 = CONVOLUTION_LOOP_for_for_for_else_and_581_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4343 = (~(CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4345 = CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4347 = CONVOLUTION_LOOP_for_for_for_else_and_579_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4349 = (~(CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4351 = CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4353 = CONVOLUTION_LOOP_for_for_for_else_and_577_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4355 = (~(CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4357 = CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4359 = CONVOLUTION_LOOP_for_for_for_else_and_575_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4361 = (~(CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4363 = CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4365 = CONVOLUTION_LOOP_for_for_for_else_and_573_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4367 = (~(CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4369 = CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4371 = CONVOLUTION_LOOP_for_for_for_else_and_571_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4373 = (~(CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4375 = CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4377 = CONVOLUTION_LOOP_for_for_for_else_and_569_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4379 = (~(CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4381 = CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4383 = CONVOLUTION_LOOP_for_for_for_else_and_567_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4385 = (~(CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4387 = CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4389 = CONVOLUTION_LOOP_for_for_for_else_and_565_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4391 = (~(CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4393 = CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4395 = CONVOLUTION_LOOP_for_for_for_else_and_563_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4397 = (~(CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4399 = CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4401 = CONVOLUTION_LOOP_for_for_for_else_and_561_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4403 = (~(CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4405 = CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4407 = CONVOLUTION_LOOP_for_for_for_else_and_559_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4409 = (~(CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4411 = CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4413 = CONVOLUTION_LOOP_for_for_for_else_and_557_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4415 = (~(CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4417 = CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4419 = CONVOLUTION_LOOP_for_for_for_else_and_555_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4421 = (~(CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4423 = CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4425 = CONVOLUTION_LOOP_for_for_for_else_and_553_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4427 = (~(CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4429 = CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4431 = CONVOLUTION_LOOP_for_for_for_else_and_551_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4433 = (~(CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4435 = CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4437 = CONVOLUTION_LOOP_for_for_for_else_and_549_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4439 = (~(CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4441 = CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4443 = CONVOLUTION_LOOP_for_for_for_else_and_547_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4445 = (~(CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4447 = CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4449 = CONVOLUTION_LOOP_for_for_for_else_and_545_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4451 = (~(CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4453 = CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4455 = CONVOLUTION_LOOP_for_for_for_else_and_543_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4457 = (~(CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4459 = CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4461 = CONVOLUTION_LOOP_for_for_for_else_and_541_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4463 = (~(CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4465 = CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4467 = CONVOLUTION_LOOP_for_for_for_else_and_539_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4469 = (~(CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4471 = CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4473 = CONVOLUTION_LOOP_for_for_for_else_and_537_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4475 = (~(CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4477 = CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4479 = CONVOLUTION_LOOP_for_for_for_else_and_535_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4481 = (~(CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4483 = CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4485 = CONVOLUTION_LOOP_for_for_for_else_and_533_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4487 = (~(CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4489 = CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4491 = CONVOLUTION_LOOP_for_for_for_else_and_531_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4493 = (~(CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4495 = CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4497 = CONVOLUTION_LOOP_for_for_for_else_and_529_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4499 = (~(CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4501 = CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4503 = CONVOLUTION_LOOP_for_for_for_else_and_527_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4505 = (~(CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4507 = CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4509 = CONVOLUTION_LOOP_for_for_for_else_and_525_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4511 = (~(CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4513 = CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4515 = CONVOLUTION_LOOP_for_for_for_else_and_523_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4517 = (~(CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4519 = CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4521 = CONVOLUTION_LOOP_for_for_for_else_and_521_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4523 = (~(CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4525 = CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4527 = CONVOLUTION_LOOP_for_for_for_else_and_519_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4529 = (~(CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4531 = CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4533 = CONVOLUTION_LOOP_for_for_for_else_and_517_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4535 = (~(CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4537 = CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4539 = CONVOLUTION_LOOP_for_for_for_else_and_515_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4541 = (~(CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4543 = CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4545 = CONVOLUTION_LOOP_for_for_for_else_and_513_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4547 = (~(CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4549 = CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4551 = CONVOLUTION_LOOP_for_for_for_else_and_512_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4553 = (~(CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4555 = CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4557 = CONVOLUTION_LOOP_for_for_for_else_and_514_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4559 = (~(CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4561 = CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4563 = CONVOLUTION_LOOP_for_for_for_else_and_516_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4565 = (~(CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4567 = CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4569 = CONVOLUTION_LOOP_for_for_for_else_and_518_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4571 = (~(CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4573 = CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4575 = CONVOLUTION_LOOP_for_for_for_else_and_520_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4577 = (~(CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4579 = CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4581 = CONVOLUTION_LOOP_for_for_for_else_and_522_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4583 = (~(CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4585 = CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4587 = CONVOLUTION_LOOP_for_for_for_else_and_524_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4589 = (~(CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4591 = CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4593 = CONVOLUTION_LOOP_for_for_for_else_and_526_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4595 = (~(CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4597 = CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4599 = CONVOLUTION_LOOP_for_for_for_else_and_528_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4601 = (~(CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4603 = CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4605 = CONVOLUTION_LOOP_for_for_for_else_and_530_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4607 = (~(CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4609 = CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4611 = CONVOLUTION_LOOP_for_for_for_else_and_532_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4613 = (~(CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4615 = CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4617 = CONVOLUTION_LOOP_for_for_for_else_and_534_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4619 = (~(CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4621 = CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4623 = CONVOLUTION_LOOP_for_for_for_else_and_536_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4625 = (~(CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4627 = CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4629 = CONVOLUTION_LOOP_for_for_for_else_and_538_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4631 = (~(CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4633 = CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4635 = CONVOLUTION_LOOP_for_for_for_else_and_540_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4637 = (~(CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4639 = CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4641 = CONVOLUTION_LOOP_for_for_for_else_and_542_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4643 = (~(CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4645 = CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4647 = CONVOLUTION_LOOP_for_for_for_else_and_544_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4649 = (~(CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4651 = CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4653 = CONVOLUTION_LOOP_for_for_for_else_and_546_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4655 = (~(CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4657 = CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4659 = CONVOLUTION_LOOP_for_for_for_else_and_548_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4661 = (~(CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4663 = CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4665 = CONVOLUTION_LOOP_for_for_for_else_and_550_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4667 = (~(CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4669 = CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4671 = CONVOLUTION_LOOP_for_for_for_else_and_552_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4673 = (~(CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4675 = CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4677 = CONVOLUTION_LOOP_for_for_for_else_and_554_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4679 = (~(CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4681 = CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4683 = CONVOLUTION_LOOP_for_for_for_else_and_556_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4685 = (~(CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4687 = CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4689 = CONVOLUTION_LOOP_for_for_for_else_and_558_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4691 = (~(CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4693 = CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4695 = CONVOLUTION_LOOP_for_for_for_else_and_560_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4697 = (~(CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4699 = CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4701 = CONVOLUTION_LOOP_for_for_for_else_and_562_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4703 = (~(CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4705 = CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4707 = CONVOLUTION_LOOP_for_for_for_else_and_564_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4709 = (~(CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4711 = CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4713 = CONVOLUTION_LOOP_for_for_for_else_and_566_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4715 = (~(CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4717 = CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4719 = CONVOLUTION_LOOP_for_for_for_else_and_568_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4721 = (~(CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4723 = CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4725 = CONVOLUTION_LOOP_for_for_for_else_and_570_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4727 = (~(CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4729 = CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4731 = CONVOLUTION_LOOP_for_for_for_else_and_572_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4733 = (~(CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4735 = CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4737 = CONVOLUTION_LOOP_for_for_for_else_and_574_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4739 = (~(CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4741 = CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4743 = CONVOLUTION_LOOP_for_for_for_else_and_576_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4745 = (~(CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4747 = CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4749 = CONVOLUTION_LOOP_for_for_for_else_and_578_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4751 = (~(CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4753 = CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4755 = CONVOLUTION_LOOP_for_for_for_else_and_580_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4757 = (~(CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4759 = CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4761 = CONVOLUTION_LOOP_for_for_for_else_and_582_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4763 = (~(CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4765 = CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4767 = CONVOLUTION_LOOP_for_for_for_else_and_584_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4769 = (~(CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4771 = CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4773 = CONVOLUTION_LOOP_for_for_for_else_and_586_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4775 = (~(CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4777 = CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4779 = CONVOLUTION_LOOP_for_for_for_else_and_588_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4781 = (~(CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4783 = CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4785 = CONVOLUTION_LOOP_for_for_for_else_and_590_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4787 = (~(CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4789 = CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4791 = CONVOLUTION_LOOP_for_for_for_else_and_592_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4793 = (~(CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4795 = CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4797 = CONVOLUTION_LOOP_for_for_for_else_and_594_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4799 = (~(CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4801 = CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4803 = CONVOLUTION_LOOP_for_for_for_else_and_596_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4805 = (~(CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4807 = CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4809 = CONVOLUTION_LOOP_for_for_for_else_and_598_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4811 = (~(CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4813 = CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4815 = CONVOLUTION_LOOP_for_for_for_else_and_600_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4817 = (~(CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4819 = CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4821 = CONVOLUTION_LOOP_for_for_for_else_and_602_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4823 = (~(CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4825 = CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4827 = CONVOLUTION_LOOP_for_for_for_else_and_604_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4829 = (~(CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4831 = CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4833 = CONVOLUTION_LOOP_for_for_for_else_and_606_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4835 = (~(CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4837 = CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4839 = CONVOLUTION_LOOP_for_for_for_else_and_608_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4841 = (~(CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4843 = CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4845 = CONVOLUTION_LOOP_for_for_for_else_and_610_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4847 = (~(CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4849 = CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4851 = CONVOLUTION_LOOP_for_for_for_else_and_612_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4853 = (~(CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4855 = CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4857 = CONVOLUTION_LOOP_for_for_for_else_and_614_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4859 = (~(CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4861 = CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4863 = CONVOLUTION_LOOP_for_for_for_else_and_616_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4865 = (~(CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4867 = CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4869 = CONVOLUTION_LOOP_for_for_for_else_and_618_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4871 = (~(CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4873 = CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4875 = CONVOLUTION_LOOP_for_for_for_else_and_620_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4877 = (~(CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4879 = CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4881 = CONVOLUTION_LOOP_for_for_for_else_and_622_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4883 = (~(CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4885 = CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4887 = CONVOLUTION_LOOP_for_for_for_else_and_624_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4889 = (~(CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4891 = CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4893 = CONVOLUTION_LOOP_for_for_for_else_and_626_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4895 = (~(CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4897 = CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4899 = CONVOLUTION_LOOP_for_for_for_else_and_628_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4901 = (~(CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4903 = CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4905 = CONVOLUTION_LOOP_for_for_for_else_and_630_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4907 = (~(CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4909 = CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4911 = CONVOLUTION_LOOP_for_for_for_else_and_632_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4913 = (~(CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4915 = CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4917 = CONVOLUTION_LOOP_for_for_for_else_and_634_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4919 = (~(CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4921 = CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4923 = CONVOLUTION_LOOP_for_for_for_else_and_636_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4925 = (~(CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4927 = CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4929 = CONVOLUTION_LOOP_for_for_for_else_and_638_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4931 = (~(CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4933 = CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4935 = CONVOLUTION_LOOP_for_for_for_else_and_640_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4937 = (~(CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4939 = CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4941 = CONVOLUTION_LOOP_for_for_for_else_and_642_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4943 = (~(CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4945 = CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4947 = CONVOLUTION_LOOP_for_for_for_else_and_644_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4949 = (~(CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4951 = CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4953 = CONVOLUTION_LOOP_for_for_for_else_and_646_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4955 = (~(CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4957 = CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4959 = CONVOLUTION_LOOP_for_for_for_else_and_648_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4961 = (~(CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4963 = CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4965 = CONVOLUTION_LOOP_for_for_for_else_and_650_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4967 = (~(CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4969 = CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4971 = CONVOLUTION_LOOP_for_for_for_else_and_652_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4973 = (~(CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4975 = CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4977 = CONVOLUTION_LOOP_for_for_for_else_and_654_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4979 = (~(CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4981 = CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4983 = CONVOLUTION_LOOP_for_for_for_else_and_656_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4985 = (~(CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4987 = CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4989 = CONVOLUTION_LOOP_for_for_for_else_and_658_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4991 = (~(CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4993 = CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4995 = CONVOLUTION_LOOP_for_for_for_else_and_660_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_4997 = (~(CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_4999 = CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5001 = CONVOLUTION_LOOP_for_for_for_else_and_662_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5003 = (~(CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5005 = CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5007 = CONVOLUTION_LOOP_for_for_for_else_and_664_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5009 = (~(CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5011 = CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5013 = CONVOLUTION_LOOP_for_for_for_else_and_666_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5015 = (~(CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5017 = CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5019 = CONVOLUTION_LOOP_for_for_for_else_and_668_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5021 = (~(CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5023 = CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5025 = CONVOLUTION_LOOP_for_for_for_else_and_670_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5027 = (~(CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5029 = CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5031 = CONVOLUTION_LOOP_for_for_for_else_and_672_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5033 = (~(CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5035 = CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5037 = CONVOLUTION_LOOP_for_for_for_else_and_674_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5039 = (~(CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5041 = CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5043 = CONVOLUTION_LOOP_for_for_for_else_and_676_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5045 = (~(CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5047 = CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5049 = CONVOLUTION_LOOP_for_for_for_else_and_678_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5051 = (~(CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5053 = CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5055 = CONVOLUTION_LOOP_for_for_for_else_and_680_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5057 = (~(CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5059 = CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5061 = CONVOLUTION_LOOP_for_for_for_else_and_682_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5063 = (~(CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5065 = CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5067 = CONVOLUTION_LOOP_for_for_for_else_and_684_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5069 = (~(CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5071 = CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5073 = CONVOLUTION_LOOP_for_for_for_else_and_686_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5075 = (~(CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5077 = CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5079 = CONVOLUTION_LOOP_for_for_for_else_and_688_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5081 = (~(CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5083 = CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5085 = CONVOLUTION_LOOP_for_for_for_else_and_690_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5087 = (~(CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5089 = CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5091 = CONVOLUTION_LOOP_for_for_for_else_and_692_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5093 = (~(CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5095 = CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5097 = CONVOLUTION_LOOP_for_for_for_else_and_694_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5099 = (~(CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5101 = CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5103 = CONVOLUTION_LOOP_for_for_for_else_and_696_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5105 = (~(CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5107 = CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5109 = CONVOLUTION_LOOP_for_for_for_else_and_698_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5111 = (~(CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5113 = CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5115 = CONVOLUTION_LOOP_for_for_for_else_and_700_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5117 = (~(CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5119 = CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5121 = CONVOLUTION_LOOP_for_for_for_else_and_702_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5123 = (~(CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5125 = CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5127 = CONVOLUTION_LOOP_for_for_for_else_and_704_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5129 = (~(CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5131 = CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5133 = CONVOLUTION_LOOP_for_for_for_else_and_706_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5135 = (~(CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5137 = CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5139 = CONVOLUTION_LOOP_for_for_for_else_and_708_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5141 = (~(CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5143 = CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5145 = CONVOLUTION_LOOP_for_for_for_else_and_710_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5147 = (~(CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5149 = CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5151 = CONVOLUTION_LOOP_for_for_for_else_and_712_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5153 = (~(CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5155 = CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5157 = CONVOLUTION_LOOP_for_for_for_else_and_714_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5159 = (~(CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5161 = CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5163 = CONVOLUTION_LOOP_for_for_for_else_and_716_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5165 = (~(CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5167 = CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5169 = CONVOLUTION_LOOP_for_for_for_else_and_718_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5171 = (~(CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5173 = CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5175 = CONVOLUTION_LOOP_for_for_for_else_and_720_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5177 = (~(CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5179 = CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5181 = CONVOLUTION_LOOP_for_for_for_else_and_722_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5183 = (~(CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5185 = CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5187 = CONVOLUTION_LOOP_for_for_for_else_and_724_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5189 = (~(CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5191 = CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5193 = CONVOLUTION_LOOP_for_for_for_else_and_726_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5195 = (~(CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5197 = CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5199 = CONVOLUTION_LOOP_for_for_for_else_and_728_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5201 = (~(CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5203 = CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5205 = CONVOLUTION_LOOP_for_for_for_else_and_730_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5207 = (~(CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5209 = CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5211 = CONVOLUTION_LOOP_for_for_for_else_and_732_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5213 = (~(CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5215 = CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5217 = CONVOLUTION_LOOP_for_for_for_else_and_734_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5219 = (~(CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5221 = CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5223 = CONVOLUTION_LOOP_for_for_for_else_and_736_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5225 = (~(CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5227 = CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5229 = CONVOLUTION_LOOP_for_for_for_else_and_738_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5231 = (~(CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5233 = CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5235 = CONVOLUTION_LOOP_for_for_for_else_and_740_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5237 = (~(CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5239 = CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5241 = CONVOLUTION_LOOP_for_for_for_else_and_742_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5243 = (~(CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5245 = CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5247 = CONVOLUTION_LOOP_for_for_for_else_and_744_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5249 = (~(CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5251 = CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5253 = CONVOLUTION_LOOP_for_for_for_else_and_746_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5255 = (~(CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5257 = CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5259 = CONVOLUTION_LOOP_for_for_for_else_and_748_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5261 = (~(CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5263 = CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5265 = CONVOLUTION_LOOP_for_for_for_else_and_750_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5267 = (~(CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5269 = CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5271 = CONVOLUTION_LOOP_for_for_for_else_and_752_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5273 = (~(CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5275 = CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5277 = CONVOLUTION_LOOP_for_for_for_else_and_754_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5279 = (~(CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5281 = CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5283 = CONVOLUTION_LOOP_for_for_for_else_and_756_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5285 = (~(CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5287 = CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5289 = CONVOLUTION_LOOP_for_for_for_else_and_758_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5291 = (~(CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5293 = CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5295 = CONVOLUTION_LOOP_for_for_for_else_and_760_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5297 = (~(CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5299 = CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5301 = CONVOLUTION_LOOP_for_for_for_else_and_762_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5303 = (~(CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5305 = CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5307 = CONVOLUTION_LOOP_for_for_for_else_and_764_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5309 = (~(CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5311 = CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5313 = CONVOLUTION_LOOP_for_for_for_else_and_766_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5315 = (~(CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5317 = CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5319 = CONVOLUTION_LOOP_for_for_for_else_and_768_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5321 = (~(CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5323 = CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5325 = CONVOLUTION_LOOP_for_for_for_else_and_770_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5327 = (~(CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5329 = CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5331 = CONVOLUTION_LOOP_for_for_for_else_and_772_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5333 = (~(CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5335 = CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5337 = CONVOLUTION_LOOP_for_for_for_else_and_774_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5339 = (~(CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5341 = CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5343 = CONVOLUTION_LOOP_for_for_for_else_and_776_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5345 = (~(CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5347 = CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5349 = CONVOLUTION_LOOP_for_for_for_else_and_778_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5351 = (~(CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5353 = CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5355 = CONVOLUTION_LOOP_for_for_for_else_and_780_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5357 = (~(CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5359 = CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5361 = CONVOLUTION_LOOP_for_for_for_else_and_782_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5363 = (~(CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5365 = CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5367 = CONVOLUTION_LOOP_for_for_for_else_and_784_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5369 = (~(CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5371 = CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5373 = CONVOLUTION_LOOP_for_for_for_else_and_786_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5375 = (~(CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5377 = CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5379 = CONVOLUTION_LOOP_for_for_for_else_and_788_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5381 = (~(CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5383 = CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5385 = CONVOLUTION_LOOP_for_for_for_else_and_790_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5387 = (~(CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5389 = CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5391 = CONVOLUTION_LOOP_for_for_for_else_and_792_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5393 = (~(CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5395 = CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5397 = CONVOLUTION_LOOP_for_for_for_else_and_794_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5399 = (~(CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5401 = CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5403 = CONVOLUTION_LOOP_for_for_for_else_and_796_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5405 = (~(CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5407 = CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5409 = CONVOLUTION_LOOP_for_for_for_else_and_798_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5411 = (~(CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5413 = CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5415 = CONVOLUTION_LOOP_for_for_for_else_and_800_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5417 = (~(CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5419 = CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5421 = CONVOLUTION_LOOP_for_for_for_else_and_802_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5423 = (~(CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5425 = CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5427 = CONVOLUTION_LOOP_for_for_for_else_and_804_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5429 = (~(CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5431 = CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5433 = CONVOLUTION_LOOP_for_for_for_else_and_806_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5435 = (~(CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5437 = CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5439 = CONVOLUTION_LOOP_for_for_for_else_and_808_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5441 = (~(CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5443 = CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5445 = CONVOLUTION_LOOP_for_for_for_else_and_810_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5447 = (~(CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5449 = CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5451 = CONVOLUTION_LOOP_for_for_for_else_and_812_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5453 = (~(CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5455 = CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5457 = CONVOLUTION_LOOP_for_for_for_else_and_814_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5459 = (~(CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5461 = CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5463 = CONVOLUTION_LOOP_for_for_for_else_and_816_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5465 = (~(CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5467 = CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5469 = CONVOLUTION_LOOP_for_for_for_else_and_818_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5471 = (~(CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5473 = CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5475 = CONVOLUTION_LOOP_for_for_for_else_and_820_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5477 = (~(CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5479 = CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5481 = CONVOLUTION_LOOP_for_for_for_else_and_822_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5483 = (~(CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5485 = CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5487 = CONVOLUTION_LOOP_for_for_for_else_and_824_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5489 = (~(CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5491 = CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5493 = CONVOLUTION_LOOP_for_for_for_else_and_826_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5495 = (~(CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5497 = CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5499 = CONVOLUTION_LOOP_for_for_for_else_and_828_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5501 = (~(CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5503 = CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5505 = CONVOLUTION_LOOP_for_for_for_else_and_830_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5507 = (~(CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5509 = CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5511 = CONVOLUTION_LOOP_for_for_for_else_and_832_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign CONVOLUTION_LOOP_for_for_for_asn_5513 = (~(CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      | CONVOLUTION_LOOP_for_for_for_unequal_tmp_1)) | ((~ CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1)
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5515 = CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      & (~ CONVOLUTION_LOOP_for_for_for_unequal_tmp_1);
  assign CONVOLUTION_LOOP_for_for_for_asn_5517 = CONVOLUTION_LOOP_for_for_for_else_and_834_ssc_sva_1
      & CONVOLUTION_LOOP_for_for_for_unequal_tmp_1;
  assign COMPUTE_LOOP_asn_44 = (~ unequal_tmp_1) & exitL_exit_COMPUTE_LOOP_sva;
  assign COMPUTE_LOOP_asn_46 = unequal_tmp_1 & exitL_exit_COMPUTE_LOOP_sva;
  assign CONVOLUTION_LOOP_for_for_for_else_CONVOLUTION_LOOP_for_for_for_else_nor_2_itm
      = ~((~((CONVOLUTION_LOOP_for_for_for_else_acc_sat_sva_1[56]) | CONVOLUTION_LOOP_for_for_for_else_and_unfl_sva_1))
      | CONVOLUTION_LOOP_for_for_for_else_nor_ovfl_sva_1);
  assign and_7_tmp = main_stage_v_1 & or_12_cse_1 & or_13_cse_1 & or_4_cse_1 & or_5_cse_1
      & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_1_cse_1 & or_2_cse_1 & or_cse_1;
  assign and_5_tmp = main_stage_v_2 & or_4_cse_1 & or_5_cse_1 & or_6_cse_1 & or_7_cse_1
      & or_8_cse_1 & or_1_cse_1 & or_2_cse_1 & or_cse_1;
  assign nor_55_cse = ~((~ operator_8_false_5_acc_itm_3_1) | CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp);
  assign or_73_cse = (~ CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp) | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)
      | (operator_8_false_1_acc_tmp[8]);
  assign and_17_nl = operator_8_false_5_acc_itm_3_1 & or_73_cse;
  assign nand_68_nl = ~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & (~(nor_55_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8]))));
  assign mux_tmp_17 = MUX_s_1_2_2(and_17_nl, nand_68_nl, operator_8_false_6_acc_itm_3_1);
  assign not_tmp_22 = ~(CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_2_CONVOLUTION_LOOP_for_for_for_if_2_nor_cse
      | (~ operator_8_false_4_acc_itm_4));
  assign or_81_nl = (~ CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp) | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)
      | (operator_8_false_1_acc_tmp[8]) | not_tmp_22;
  assign mux_34_nl = MUX_s_1_2_2(not_tmp_22, or_81_nl, operator_8_false_5_acc_itm_3_1);
  assign nand_69_nl = ~(CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp & (~(nor_55_cse
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8])
      | not_tmp_22)));
  assign mux_35_cse = MUX_s_1_2_2(mux_34_nl, nand_69_nl, operator_8_false_6_acc_itm_3_1);
  assign or_tmp_46 = (CONVOLUTION_LOOP_for_for_if_or_cse & operator_8_false_3_acc_itm_4_1)
      | mux_35_cse;
  assign nor_40_cse = ~((~((operator_8_false_3_acc_tmp[8:5]!=4'b0000) | (~ CONVOLUTION_LOOP_for_if_equal_tmp)))
      | (CONVOLUTION_LOOP_for_acc_tmp[5]));
  assign nand_tmp_7 = nor_40_cse | or_tmp_46;
  assign or_87_nl = CONVOLUTION_LOOP_if_CONVOLUTION_LOOP_if_nand_tmp | (operator_8_false_7_acc_tmp[8])
      | nand_tmp_7;
  assign mux_tmp_21 = MUX_s_1_2_2(or_87_nl, nand_tmp_7, CONVOLUTION_LOOP_acc_tmp[5]);
  assign and_dcpl_7 = and_9_tmp & COMPUTE_LOOP_asn_itm;
  assign and_dcpl_11 = exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_2 & and_5_tmp;
  assign and_dcpl_17 = ~(exitL_exit_COMPUTE_LOOP_sva | exit_COMPUTE_LOOP_lpi_1_dfm_2);
  assign and_dcpl_19 = (~((~(and_dcpl_17 & (~ exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1)))
      & and_9_tmp)) & and_235_cse;
  assign or_dcpl_14 = plm_outputs_rsci_bawt | (~ CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3)
      | (~ exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_3);
  assign or_dcpl_15 = (~ exit_COMPUTE_LOOP_lpi_1_dfm_2_st_4) | done_rsci_bawt;
  assign or_dcpl_16 = or_dcpl_15 | (~ main_stage_v_4);
  assign and_dcpl_28 = or_dcpl_16 & (plm_outputs_rsc_rls_obj_bawt | (~ exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_3));
  assign and_dcpl_29 = and_dcpl_28 & or_dcpl_14;
  assign and_dcpl_32 = exit_COMPUTE_LOOP_lpi_1_dfm_2_st_4 & done_rsci_bawt & main_stage_v_4;
  assign and_dcpl_36 = (and_10_cse | and_11_cse | (~ main_stage_v_3) | (~ exit_COMPUTE_LOOP_lpi_1_dfm_2_st_3))
      & and_dcpl_32;
  assign or_dcpl_22 = ~(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_2 &
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2
      & and_5_tmp);
  assign or_dcpl_31 = ~(exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_2 &
      and_5_tmp);
  assign and_dcpl_57 = (~((~((~ (operator_8_false_1_acc_tmp[8])) & CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp
      & CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp)) & operator_8_false_6_acc_itm_3_1))
      & and_9_tmp;
  assign or_dcpl_34 = (operator_8_false_1_acc_tmp[8]) | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp)
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp);
  assign and_dcpl_59 = or_dcpl_34 & operator_8_false_6_acc_itm_3_1 & and_9_tmp;
  assign or_dcpl_39 = ~(exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0 & and_9_tmp);
  assign or_dcpl_40 = nor_40_cse | mux_tmp_17 | not_tmp_22;
  assign and_dcpl_66 = or_dcpl_34 & operator_8_false_6_acc_itm_3_1;
  assign and_dcpl_72 = (~ or_dcpl_40) & exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0
      & and_9_tmp;
  assign and_dcpl_73 = nand_tmp_7 & and_9_tmp;
  assign and_dcpl_84 = (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0)
      & and_dcpl_17 & (~(exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1 | exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3))
      & (~(exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3 | exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2));
  assign or_tmp_98 = (mux_tmp_21 | (~((exit_COMPUTE_LOOP_sva_2_mx0w0 | (COMPUTE_LOOP_acc_tmp[4]))
      & and_9_tmp))) & and_dcpl_7 & (fsm_output[1]);
  assign and_113_cse = COMPUTE_LOOP_COMPUTE_LOOP_or_tmp & and_9_tmp & (fsm_output[1]);
  assign or_tmp_108 = and_7_tmp & (fsm_output[1]);
  assign or_tmp_109 = and_5_tmp & (fsm_output[1]);
  assign or_tmp_111 = (~ and_7_tmp) | (fsm_output[0]);
  assign plm_outputs_rsc_req_obj_iswt0_mx0c1 = (~(and_7_tmp & exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_1))
      & and_dcpl_11;
  assign main_stage_v_3_mx0c1 = and_dcpl_29 & main_stage_v_3 & (~ and_5_tmp);
  assign main_stage_v_4_mx0c1 = (and_10_cse | and_11_cse | (~ main_stage_v_3)) &
      or_dcpl_15 & main_stage_v_4;
  assign main_stage_v_2_mx0c1 = (~ and_7_tmp) & and_5_tmp & (fsm_output[1]);
  assign main_stage_v_1_mx0c1 = and_7_tmp & (~ and_9_tmp) & (fsm_output[1]);
  assign CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1
      = mux_tmp_17 & and_9_tmp & (fsm_output[1]);
  assign nl_operator_8_false_6_acc_nl = ({1'b1 , CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2})
      + 4'b0001;
  assign operator_8_false_6_acc_nl = nl_operator_8_false_6_acc_nl[3:0];
  assign operator_8_false_6_acc_itm_3_1 = readslicef_4_1_3(operator_8_false_6_acc_nl);
  assign plm_inputs_rsci_radr_d = CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff;
  assign plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign plm_filters_rsci_radr_d = CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff;
  assign plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign plm_outputs_rsci_d_d = {CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff , CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff
      , CONVOLUTION_LOOP_for_for_for_if_1_mux_rmff};
  assign plm_outputs_rsci_wadr_d = CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff;
  assign plm_outputs_rsci_we_d_pff = plm_outputs_rsci_we_d_iff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (((~ mux_37_nl) & and_9_tmp) | (fsm_output[0]) | or_tmp_98)
        ) begin
      reg_conf_info_rsci_iswt0_cse <= ~ or_tmp_98;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exitL_exit_COMPUTE_LOOP_sva <= 1'b1;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_1 <= 1'b0;
      exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1 <= 14'b00000000000000;
      CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1 <= 16'b0000000000000000;
      exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      exit_COMPUTE_LOOP_lpi_1_dfm_2 <= 1'b0;
      exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3 <= 1'b0;
      exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3 <= 1'b0;
      exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2 <= 1'b0;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( COMPUTE_LOOP_and_cse ) begin
      exitL_exit_COMPUTE_LOOP_sva <= exit_COMPUTE_LOOP_lpi_1_dfm_2_mx0w0;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_1 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_mx0w0;
      exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1 <= exit_CONVOLUTION_LOOP_lpi_1_dfm_3_mx0w0;
      CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1 <= nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1[13:0];
      CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1 <= nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1[15:0];
      exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_1 <= COMPUTE_LOOP_COMPUTE_LOOP_or_tmp;
      exit_COMPUTE_LOOP_lpi_1_dfm_2 <= exit_COMPUTE_LOOP_lpi_1_dfm_2_mx0w0;
      exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3 <= exit_CONVOLUTION_LOOP_for_lpi_1_dfm_3_mx0w0;
      exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3 <= exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_3_mx0w0;
      exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2 <= exit_CONVOLUTION_LOOP_for_for_for_lpi_1_dfm_2_mx0w0;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsc_req_obj_iswt0 <= 1'b0;
    end
    else if ( core_wen & (and_235_cse | plm_outputs_rsc_req_obj_iswt0_mx0c1) ) begin
      plm_outputs_rsc_req_obj_iswt0 <= ~ plm_outputs_rsc_req_obj_iswt0_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_inputs_rsc_req_obj_iswt0 <= 1'b0;
    end
    else if ( core_wen & (and_113_cse | ((exit_COMPUTE_LOOP_lpi_1_dfm_2 | exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1)
        & (~ exitL_exit_COMPUTE_LOOP_sva) & and_9_tmp) | and_dcpl_19) ) begin
      plm_inputs_rsc_req_obj_iswt0 <= ~ and_dcpl_19;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_filters_rsc_req_obj_iswt0 <= 1'b0;
    end
    else if ( core_wen & (and_113_cse | and_dcpl_19) ) begin
      plm_filters_rsc_req_obj_iswt0 <= ~ and_dcpl_19;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_filters_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_plm_filters_rsc_rls_obj_oswt_cse <= 1'b0;
      reg_plm_outputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= 1'b0;
      reg_plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
      plm_outputs_rsci_wadr_d_reg <= 14'b00000000000000;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5 <=
          1'b0;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4 <=
          30'b000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3 <=
          1'b0;
      plm_filters_rsci_radr_d_reg <= 16'b0000000000000000;
      plm_inputs_rsci_radr_d_reg <= 14'b00000000000000;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1 <= 1'b0;
      lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1 <= 1'b0;
      conf_info_crt_lpi_1_dfm_231_224 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_71_64 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_135_128 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_103_96 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_7_0 <= 8'b00000000;
      n_w_in_acc_psp_lpi_1_dfm <= 7'b0000000;
      conf_info_crt_lpi_1_dfm_192 <= 1'b0;
      n_h_in_acc_psp_lpi_1_dfm <= 7'b0000000;
      conf_info_crt_lpi_1_dfm_160 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_plm_filters_rsc_rls_obj_ld_core_psct_cse <= and_7_tmp & exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1;
      reg_plm_filters_rsc_rls_obj_oswt_cse <= and_34_rmff;
      reg_plm_outputs_rsci_writeA_w_ram_ir_internal_WMASK_B_d_core_psct_cse <= and_50_rmff;
      reg_plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= or_tmp_108;
      plm_outputs_rsci_wadr_d_reg <= CONVOLUTION_LOOP_for_for_for_index_out_mux_rmff;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_5 <=
          CONVOLUTION_LOOP_for_for_for_if_1_mux_rmff;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_4 <=
          CONVOLUTION_LOOP_for_for_for_if_1_mux_3_rmff;
      CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_3 <=
          CONVOLUTION_LOOP_for_for_for_if_1_mux_4_rmff;
      plm_filters_rsci_radr_d_reg <= CONVOLUTION_LOOP_for_for_for_for_for_mux_rmff;
      plm_inputs_rsci_radr_d_reg <= CONVOLUTION_LOOP_for_for_for_for_for_mux_1_rmff;
      exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1 <= exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0;
      lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1 <= lfst_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_mx0;
      conf_info_crt_lpi_1_dfm_231_224 <= conf_info_crt_lpi_1_dfm_231_224_mx0;
      conf_info_crt_lpi_1_dfm_71_64 <= conf_info_crt_lpi_1_dfm_71_64_mx0;
      conf_info_crt_lpi_1_dfm_135_128 <= conf_info_crt_lpi_1_dfm_135_128_mx0;
      conf_info_crt_lpi_1_dfm_103_96 <= conf_info_crt_lpi_1_dfm_103_96_mx0;
      conf_info_crt_lpi_1_dfm_7_0 <= conf_info_crt_lpi_1_dfm_7_0_mx0;
      n_w_in_acc_psp_lpi_1_dfm <= n_w_in_acc_psp_lpi_1_dfm_mx0;
      conf_info_crt_lpi_1_dfm_192 <= conf_info_crt_lpi_1_dfm_192_mx0;
      n_h_in_acc_psp_lpi_1_dfm <= n_h_in_acc_psp_lpi_1_dfm_mx0;
      conf_info_crt_lpi_1_dfm_160 <= conf_info_crt_lpi_1_dfm_160_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_done_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & main_stage_v_3 & exit_COMPUTE_LOOP_lpi_1_dfm_2_st_3)
        | and_dcpl_36) ) begin
      reg_done_rsci_ivld_core_psct_cse <= ~ and_dcpl_36;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_LOOP_asn_itm <= 1'b1;
    end
    else if ( core_wen & and_131_cse ) begin
      COMPUTE_LOOP_asn_itm <= exit_COMPUTE_LOOP_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_109 | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
          <= 1'b0;
      exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_3 <= 1'b0;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_3 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1 <= 45'b000000000000000000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_acc_46_sva_1 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_if_1_and_cse ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_3
          <= CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2;
      exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_3 <= exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_2;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_3 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_2;
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1 <= CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0;
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1 <= CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0;
      CONVOLUTION_LOOP_for_for_for_acc_46_sva_1 <= CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_2_st_3 <= 1'b0;
    end
    else if ( core_wen & and_5_tmp ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_2_st_3 <= exit_COMPUTE_LOOP_lpi_1_dfm_2_st_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_29 & main_stage_v_3) | main_stage_v_4_mx0c1)
        ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_2_st_4 <= 1'b0;
    end
    else if ( core_wen & (~((exit_COMPUTE_LOOP_lpi_1_dfm_2_st_4 & (~ done_rsci_bawt)
        & main_stage_v_4) | and_11_cse | and_10_cse | (~ main_stage_v_3))) ) begin
      exit_COMPUTE_LOOP_lpi_1_dfm_2_st_4 <= exit_COMPUTE_LOOP_lpi_1_dfm_2_st_3;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_108 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_2 <= 11'b00000000000;
      COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_2 <= 1'b0;
      COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_2 <= 45'b000000000000000000000000000000000000000000000;
      COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_2 <= 11'b00000000000;
    end
    else if ( COMPUTE_LOOP_buf_acc_data_and_cse ) begin
      COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_1_mx0;
      COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_3;
      COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_2 <= COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_3;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0 <= 1'b0;
      reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse <= 5'b00000;
      reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_else_mux_itm_1 <= 11'b00000000000;
      CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1 <= 45'b000000000000000000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2 <= 14'b00000000000000;
      CONVOLUTION_LOOP_for_for_for_unequal_tmp_1 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_j_and_cse ) begin
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_2_0 <= CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1_0;
      reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_7_3_cse <= CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3;
      reg_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_2_2_0_cse <= CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0;
      CONVOLUTION_LOOP_for_for_for_else_mux_itm_1 <= MUX_v_11_324_2(CONVOLUTION_LOOP_for_for_for_for_mux_12_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_24_nl, CONVOLUTION_LOOP_for_for_for_for_mux_36_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_48_nl, CONVOLUTION_LOOP_for_for_for_for_mux_60_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_72_nl, CONVOLUTION_LOOP_for_for_for_for_mux_84_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_96_nl, CONVOLUTION_LOOP_for_for_for_for_mux_108_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_120_nl, CONVOLUTION_LOOP_for_for_for_for_mux_132_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_144_nl, CONVOLUTION_LOOP_for_for_for_for_mux_156_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_168_nl, CONVOLUTION_LOOP_for_for_for_for_mux_180_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_192_nl, CONVOLUTION_LOOP_for_for_for_for_mux_204_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_216_nl, CONVOLUTION_LOOP_for_for_for_for_mux_228_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_240_nl, CONVOLUTION_LOOP_for_for_for_for_mux_252_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_264_nl, CONVOLUTION_LOOP_for_for_for_for_mux_276_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_288_nl, CONVOLUTION_LOOP_for_for_for_for_mux_300_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_312_nl, CONVOLUTION_LOOP_for_for_for_for_mux_324_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_336_nl, CONVOLUTION_LOOP_for_for_for_for_mux_348_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_360_nl, CONVOLUTION_LOOP_for_for_for_for_mux_372_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_384_nl, CONVOLUTION_LOOP_for_for_for_for_mux_396_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_408_nl, CONVOLUTION_LOOP_for_for_for_for_mux_420_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_432_nl, CONVOLUTION_LOOP_for_for_for_for_mux_444_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_456_nl, CONVOLUTION_LOOP_for_for_for_for_mux_468_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_480_nl, CONVOLUTION_LOOP_for_for_for_for_mux_492_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_504_nl, CONVOLUTION_LOOP_for_for_for_for_mux_516_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_528_nl, CONVOLUTION_LOOP_for_for_for_for_mux_540_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_552_nl, CONVOLUTION_LOOP_for_for_for_for_mux_564_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_576_nl, CONVOLUTION_LOOP_for_for_for_for_mux_588_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_600_nl, CONVOLUTION_LOOP_for_for_for_for_mux_612_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_624_nl, CONVOLUTION_LOOP_for_for_for_for_mux_636_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_648_nl, CONVOLUTION_LOOP_for_for_for_for_mux_660_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_672_nl, CONVOLUTION_LOOP_for_for_for_for_mux_684_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_696_nl, CONVOLUTION_LOOP_for_for_for_for_mux_708_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_720_nl, CONVOLUTION_LOOP_for_for_for_for_mux_732_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_744_nl, CONVOLUTION_LOOP_for_for_for_for_mux_756_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_768_nl, CONVOLUTION_LOOP_for_for_for_for_mux_780_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_792_nl, CONVOLUTION_LOOP_for_for_for_for_mux_804_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_816_nl, CONVOLUTION_LOOP_for_for_for_for_mux_828_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_840_nl, CONVOLUTION_LOOP_for_for_for_for_mux_852_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_864_nl, CONVOLUTION_LOOP_for_for_for_for_mux_876_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_888_nl, CONVOLUTION_LOOP_for_for_for_for_mux_900_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_912_nl, CONVOLUTION_LOOP_for_for_for_for_mux_924_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_936_nl, CONVOLUTION_LOOP_for_for_for_for_mux_948_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_960_nl, CONVOLUTION_LOOP_for_for_for_for_mux_972_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_984_nl, CONVOLUTION_LOOP_for_for_for_for_mux_996_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1008_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1020_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1032_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1044_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1056_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1068_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1080_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1092_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1104_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1116_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1128_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1140_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1152_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1164_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1176_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1188_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1200_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1212_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1224_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1236_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1248_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1260_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1272_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1284_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1296_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1308_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1320_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1332_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1344_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1356_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1368_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1380_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1392_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1404_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1416_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1428_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1440_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1452_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1464_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1476_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1488_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1500_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1512_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1524_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1536_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1548_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1560_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1572_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1584_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1596_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1608_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1620_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1632_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1644_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1656_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1668_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1680_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1692_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1704_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1716_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1728_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1740_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1752_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1764_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1776_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1788_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1800_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1812_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1824_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1836_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1848_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1860_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1872_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1884_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1896_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1908_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1920_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1932_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1944_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1938_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1926_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1914_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1902_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1890_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1878_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1866_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1854_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1842_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1830_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1818_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1806_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1794_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1782_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1770_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1758_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1746_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1734_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1722_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1710_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1698_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1686_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1674_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1662_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1650_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1638_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1626_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1614_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1602_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1590_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1578_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1566_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1554_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1542_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1530_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1518_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1506_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1494_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1482_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1470_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1458_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1446_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1434_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1422_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1410_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1398_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1386_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1374_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1362_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1350_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1338_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1326_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1314_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1302_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1290_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1278_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1266_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1254_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1242_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1230_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1218_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1206_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1194_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1182_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1170_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1158_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1146_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1134_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1122_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1110_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1098_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1086_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1074_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1062_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1050_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1038_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1026_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1014_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1002_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_990_nl, CONVOLUTION_LOOP_for_for_for_for_mux_978_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_966_nl, CONVOLUTION_LOOP_for_for_for_for_mux_954_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_942_nl, CONVOLUTION_LOOP_for_for_for_for_mux_930_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_918_nl, CONVOLUTION_LOOP_for_for_for_for_mux_906_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_894_nl, CONVOLUTION_LOOP_for_for_for_for_mux_882_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_870_nl, CONVOLUTION_LOOP_for_for_for_for_mux_858_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_846_nl, CONVOLUTION_LOOP_for_for_for_for_mux_834_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_822_nl, CONVOLUTION_LOOP_for_for_for_for_mux_810_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_798_nl, CONVOLUTION_LOOP_for_for_for_for_mux_786_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_774_nl, CONVOLUTION_LOOP_for_for_for_for_mux_762_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_750_nl, CONVOLUTION_LOOP_for_for_for_for_mux_738_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_726_nl, CONVOLUTION_LOOP_for_for_for_for_mux_714_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_702_nl, CONVOLUTION_LOOP_for_for_for_for_mux_690_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_678_nl, CONVOLUTION_LOOP_for_for_for_for_mux_666_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_654_nl, CONVOLUTION_LOOP_for_for_for_for_mux_642_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_630_nl, CONVOLUTION_LOOP_for_for_for_for_mux_618_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_606_nl, CONVOLUTION_LOOP_for_for_for_for_mux_594_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_582_nl, CONVOLUTION_LOOP_for_for_for_for_mux_570_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_558_nl, CONVOLUTION_LOOP_for_for_for_for_mux_546_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_534_nl, CONVOLUTION_LOOP_for_for_for_for_mux_522_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_510_nl, CONVOLUTION_LOOP_for_for_for_for_mux_498_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_486_nl, CONVOLUTION_LOOP_for_for_for_for_mux_474_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_462_nl, CONVOLUTION_LOOP_for_for_for_for_mux_450_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_438_nl, CONVOLUTION_LOOP_for_for_for_for_mux_426_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_414_nl, CONVOLUTION_LOOP_for_for_for_for_mux_402_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_390_nl, CONVOLUTION_LOOP_for_for_for_for_mux_378_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_366_nl, CONVOLUTION_LOOP_for_for_for_for_mux_354_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_342_nl, CONVOLUTION_LOOP_for_for_for_for_mux_330_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_318_nl, CONVOLUTION_LOOP_for_for_for_for_mux_306_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_294_nl, CONVOLUTION_LOOP_for_for_for_for_mux_282_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_270_nl, CONVOLUTION_LOOP_for_for_for_for_mux_258_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_246_nl, CONVOLUTION_LOOP_for_for_for_for_mux_234_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_222_nl, CONVOLUTION_LOOP_for_for_for_for_mux_210_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_198_nl, CONVOLUTION_LOOP_for_for_for_for_mux_186_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_174_nl, CONVOLUTION_LOOP_for_for_for_for_mux_162_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_150_nl, CONVOLUTION_LOOP_for_for_for_for_mux_138_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_126_nl, CONVOLUTION_LOOP_for_for_for_for_mux_114_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_102_nl, CONVOLUTION_LOOP_for_for_for_for_mux_90_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_78_nl, CONVOLUTION_LOOP_for_for_for_for_mux_66_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_54_nl, CONVOLUTION_LOOP_for_for_for_for_mux_42_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_30_nl, CONVOLUTION_LOOP_for_for_for_for_mux_18_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_6_nl, {CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3
          , CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1_0});
      CONVOLUTION_LOOP_for_for_for_else_mux_972_itm_1 <= MUX_v_45_324_2(CONVOLUTION_LOOP_for_for_for_for_mux_10_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_22_nl, CONVOLUTION_LOOP_for_for_for_for_mux_34_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_46_nl, CONVOLUTION_LOOP_for_for_for_for_mux_58_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_70_nl, CONVOLUTION_LOOP_for_for_for_for_mux_82_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_94_nl, CONVOLUTION_LOOP_for_for_for_for_mux_106_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_118_nl, CONVOLUTION_LOOP_for_for_for_for_mux_130_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_142_nl, CONVOLUTION_LOOP_for_for_for_for_mux_154_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_166_nl, CONVOLUTION_LOOP_for_for_for_for_mux_178_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_190_nl, CONVOLUTION_LOOP_for_for_for_for_mux_202_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_214_nl, CONVOLUTION_LOOP_for_for_for_for_mux_226_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_238_nl, CONVOLUTION_LOOP_for_for_for_for_mux_250_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_262_nl, CONVOLUTION_LOOP_for_for_for_for_mux_274_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_286_nl, CONVOLUTION_LOOP_for_for_for_for_mux_298_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_310_nl, CONVOLUTION_LOOP_for_for_for_for_mux_322_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_334_nl, CONVOLUTION_LOOP_for_for_for_for_mux_346_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_358_nl, CONVOLUTION_LOOP_for_for_for_for_mux_370_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_382_nl, CONVOLUTION_LOOP_for_for_for_for_mux_394_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_406_nl, CONVOLUTION_LOOP_for_for_for_for_mux_418_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_430_nl, CONVOLUTION_LOOP_for_for_for_for_mux_442_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_454_nl, CONVOLUTION_LOOP_for_for_for_for_mux_466_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_478_nl, CONVOLUTION_LOOP_for_for_for_for_mux_490_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_502_nl, CONVOLUTION_LOOP_for_for_for_for_mux_514_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_526_nl, CONVOLUTION_LOOP_for_for_for_for_mux_538_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_550_nl, CONVOLUTION_LOOP_for_for_for_for_mux_562_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_574_nl, CONVOLUTION_LOOP_for_for_for_for_mux_586_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_598_nl, CONVOLUTION_LOOP_for_for_for_for_mux_610_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_622_nl, CONVOLUTION_LOOP_for_for_for_for_mux_634_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_646_nl, CONVOLUTION_LOOP_for_for_for_for_mux_658_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_670_nl, CONVOLUTION_LOOP_for_for_for_for_mux_682_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_694_nl, CONVOLUTION_LOOP_for_for_for_for_mux_706_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_718_nl, CONVOLUTION_LOOP_for_for_for_for_mux_730_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_742_nl, CONVOLUTION_LOOP_for_for_for_for_mux_754_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_766_nl, CONVOLUTION_LOOP_for_for_for_for_mux_778_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_790_nl, CONVOLUTION_LOOP_for_for_for_for_mux_802_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_814_nl, CONVOLUTION_LOOP_for_for_for_for_mux_826_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_838_nl, CONVOLUTION_LOOP_for_for_for_for_mux_850_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_862_nl, CONVOLUTION_LOOP_for_for_for_for_mux_874_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_886_nl, CONVOLUTION_LOOP_for_for_for_for_mux_898_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_910_nl, CONVOLUTION_LOOP_for_for_for_for_mux_922_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_934_nl, CONVOLUTION_LOOP_for_for_for_for_mux_946_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_958_nl, CONVOLUTION_LOOP_for_for_for_for_mux_970_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_982_nl, CONVOLUTION_LOOP_for_for_for_for_mux_994_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1006_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1018_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1030_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1042_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1054_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1066_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1078_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1090_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1102_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1114_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1126_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1138_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1150_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1162_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1174_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1186_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1198_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1210_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1222_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1234_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1246_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1258_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1270_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1282_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1294_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1306_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1318_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1330_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1342_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1354_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1366_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1378_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1390_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1402_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1414_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1426_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1438_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1450_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1462_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1474_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1486_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1498_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1510_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1522_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1534_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1546_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1558_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1570_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1582_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1594_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1606_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1618_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1630_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1642_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1654_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1666_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1678_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1690_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1702_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1714_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1726_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1738_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1750_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1762_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1774_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1786_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1798_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1810_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1822_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1834_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1846_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1858_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1870_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1882_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1894_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1906_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1918_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1930_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1942_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1936_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1924_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1912_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1900_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1888_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1876_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1864_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1852_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1840_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1828_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1816_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1804_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1792_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1780_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1768_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1756_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1744_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1732_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1720_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1708_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1696_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1684_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1672_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1660_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1648_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1636_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1624_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1612_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1600_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1588_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1576_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1564_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1552_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1540_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1528_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1516_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1504_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1492_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1480_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1468_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1456_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1444_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1432_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1420_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1408_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1396_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1384_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1372_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1360_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1348_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1336_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1324_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1312_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1300_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1288_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1276_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1264_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1252_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1240_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1228_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1216_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1204_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1192_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1180_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1168_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1156_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1144_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1132_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1120_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1108_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1096_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1084_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1072_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1060_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1048_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1036_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1024_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1012_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1000_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_988_nl, CONVOLUTION_LOOP_for_for_for_for_mux_976_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_964_nl, CONVOLUTION_LOOP_for_for_for_for_mux_952_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_940_nl, CONVOLUTION_LOOP_for_for_for_for_mux_928_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_916_nl, CONVOLUTION_LOOP_for_for_for_for_mux_904_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_892_nl, CONVOLUTION_LOOP_for_for_for_for_mux_880_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_868_nl, CONVOLUTION_LOOP_for_for_for_for_mux_856_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_844_nl, CONVOLUTION_LOOP_for_for_for_for_mux_832_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_820_nl, CONVOLUTION_LOOP_for_for_for_for_mux_808_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_796_nl, CONVOLUTION_LOOP_for_for_for_for_mux_784_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_772_nl, CONVOLUTION_LOOP_for_for_for_for_mux_760_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_748_nl, CONVOLUTION_LOOP_for_for_for_for_mux_736_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_724_nl, CONVOLUTION_LOOP_for_for_for_for_mux_712_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_700_nl, CONVOLUTION_LOOP_for_for_for_for_mux_688_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_676_nl, CONVOLUTION_LOOP_for_for_for_for_mux_664_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_652_nl, CONVOLUTION_LOOP_for_for_for_for_mux_640_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_628_nl, CONVOLUTION_LOOP_for_for_for_for_mux_616_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_604_nl, CONVOLUTION_LOOP_for_for_for_for_mux_592_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_580_nl, CONVOLUTION_LOOP_for_for_for_for_mux_568_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_556_nl, CONVOLUTION_LOOP_for_for_for_for_mux_544_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_532_nl, CONVOLUTION_LOOP_for_for_for_for_mux_520_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_508_nl, CONVOLUTION_LOOP_for_for_for_for_mux_496_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_484_nl, CONVOLUTION_LOOP_for_for_for_for_mux_472_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_460_nl, CONVOLUTION_LOOP_for_for_for_for_mux_448_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_436_nl, CONVOLUTION_LOOP_for_for_for_for_mux_424_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_412_nl, CONVOLUTION_LOOP_for_for_for_for_mux_400_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_388_nl, CONVOLUTION_LOOP_for_for_for_for_mux_376_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_364_nl, CONVOLUTION_LOOP_for_for_for_for_mux_352_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_340_nl, CONVOLUTION_LOOP_for_for_for_for_mux_328_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_316_nl, CONVOLUTION_LOOP_for_for_for_for_mux_304_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_292_nl, CONVOLUTION_LOOP_for_for_for_for_mux_280_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_268_nl, CONVOLUTION_LOOP_for_for_for_for_mux_256_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_244_nl, CONVOLUTION_LOOP_for_for_for_for_mux_232_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_220_nl, CONVOLUTION_LOOP_for_for_for_for_mux_208_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_196_nl, CONVOLUTION_LOOP_for_for_for_for_mux_184_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_172_nl, CONVOLUTION_LOOP_for_for_for_for_mux_160_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_148_nl, CONVOLUTION_LOOP_for_for_for_for_mux_136_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_124_nl, CONVOLUTION_LOOP_for_for_for_for_mux_112_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_100_nl, CONVOLUTION_LOOP_for_for_for_for_mux_88_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_76_nl, CONVOLUTION_LOOP_for_for_for_for_mux_64_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_52_nl, CONVOLUTION_LOOP_for_for_for_for_mux_40_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_28_nl, CONVOLUTION_LOOP_for_for_for_for_mux_16_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_4_nl, {CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3
          , CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1_0});
      CONVOLUTION_LOOP_for_for_for_else_mux_973_itm_1 <= MUX_s_1_324_2(CONVOLUTION_LOOP_for_for_for_for_mux_8_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_20_nl, CONVOLUTION_LOOP_for_for_for_for_mux_32_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_44_nl, CONVOLUTION_LOOP_for_for_for_for_mux_56_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_68_nl, CONVOLUTION_LOOP_for_for_for_for_mux_80_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_92_nl, CONVOLUTION_LOOP_for_for_for_for_mux_104_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_116_nl, CONVOLUTION_LOOP_for_for_for_for_mux_128_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_140_nl, CONVOLUTION_LOOP_for_for_for_for_mux_152_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_164_nl, CONVOLUTION_LOOP_for_for_for_for_mux_176_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_188_nl, CONVOLUTION_LOOP_for_for_for_for_mux_200_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_212_nl, CONVOLUTION_LOOP_for_for_for_for_mux_224_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_236_nl, CONVOLUTION_LOOP_for_for_for_for_mux_248_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_260_nl, CONVOLUTION_LOOP_for_for_for_for_mux_272_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_284_nl, CONVOLUTION_LOOP_for_for_for_for_mux_296_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_308_nl, CONVOLUTION_LOOP_for_for_for_for_mux_320_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_332_nl, CONVOLUTION_LOOP_for_for_for_for_mux_344_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_356_nl, CONVOLUTION_LOOP_for_for_for_for_mux_368_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_380_nl, CONVOLUTION_LOOP_for_for_for_for_mux_392_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_404_nl, CONVOLUTION_LOOP_for_for_for_for_mux_416_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_428_nl, CONVOLUTION_LOOP_for_for_for_for_mux_440_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_452_nl, CONVOLUTION_LOOP_for_for_for_for_mux_464_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_476_nl, CONVOLUTION_LOOP_for_for_for_for_mux_488_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_500_nl, CONVOLUTION_LOOP_for_for_for_for_mux_512_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_524_nl, CONVOLUTION_LOOP_for_for_for_for_mux_536_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_548_nl, CONVOLUTION_LOOP_for_for_for_for_mux_560_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_572_nl, CONVOLUTION_LOOP_for_for_for_for_mux_584_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_596_nl, CONVOLUTION_LOOP_for_for_for_for_mux_608_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_620_nl, CONVOLUTION_LOOP_for_for_for_for_mux_632_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_644_nl, CONVOLUTION_LOOP_for_for_for_for_mux_656_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_668_nl, CONVOLUTION_LOOP_for_for_for_for_mux_680_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_692_nl, CONVOLUTION_LOOP_for_for_for_for_mux_704_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_716_nl, CONVOLUTION_LOOP_for_for_for_for_mux_728_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_740_nl, CONVOLUTION_LOOP_for_for_for_for_mux_752_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_764_nl, CONVOLUTION_LOOP_for_for_for_for_mux_776_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_788_nl, CONVOLUTION_LOOP_for_for_for_for_mux_800_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_812_nl, CONVOLUTION_LOOP_for_for_for_for_mux_824_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_836_nl, CONVOLUTION_LOOP_for_for_for_for_mux_848_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_860_nl, CONVOLUTION_LOOP_for_for_for_for_mux_872_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_884_nl, CONVOLUTION_LOOP_for_for_for_for_mux_896_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_908_nl, CONVOLUTION_LOOP_for_for_for_for_mux_920_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_932_nl, CONVOLUTION_LOOP_for_for_for_for_mux_944_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_956_nl, CONVOLUTION_LOOP_for_for_for_for_mux_968_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_980_nl, CONVOLUTION_LOOP_for_for_for_for_mux_992_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1004_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1016_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1028_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1040_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1052_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1064_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1076_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1088_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1100_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1112_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1124_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1136_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1148_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1160_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1172_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1184_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1196_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1208_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1220_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1232_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1244_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1256_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1268_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1280_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1292_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1304_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1316_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1328_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1340_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1352_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1364_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1376_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1388_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1400_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1412_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1424_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1436_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1448_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1460_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1472_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1484_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1496_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1508_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1520_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1532_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1544_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1556_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1568_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1580_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1592_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1604_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1616_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1628_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1640_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1652_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1664_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1676_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1688_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1700_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1712_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1724_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1736_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1748_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1760_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1772_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1784_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1796_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1808_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1820_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1832_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1844_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1856_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1868_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1880_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1892_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1904_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1916_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1928_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1940_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1934_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1922_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1910_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1898_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1886_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1874_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1862_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1850_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1838_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1826_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1814_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1802_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1790_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1778_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1766_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1754_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1742_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1730_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1718_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1706_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1694_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1682_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1670_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1658_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1646_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1634_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1622_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1610_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1598_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1586_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1574_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1562_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1550_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1538_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1526_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1514_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1502_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1490_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1478_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1466_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1454_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1442_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1430_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1418_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1406_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1394_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1382_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1370_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1358_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1346_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1334_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1322_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1310_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1298_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1286_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1274_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1262_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1250_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1238_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1226_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1214_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1202_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1190_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1178_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1166_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1154_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1142_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1130_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1118_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1106_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1094_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1082_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1070_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1058_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1046_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1034_nl, CONVOLUTION_LOOP_for_for_for_for_mux_1022_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_1010_nl, CONVOLUTION_LOOP_for_for_for_for_mux_998_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_986_nl, CONVOLUTION_LOOP_for_for_for_for_mux_974_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_962_nl, CONVOLUTION_LOOP_for_for_for_for_mux_950_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_938_nl, CONVOLUTION_LOOP_for_for_for_for_mux_926_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_914_nl, CONVOLUTION_LOOP_for_for_for_for_mux_902_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_890_nl, CONVOLUTION_LOOP_for_for_for_for_mux_878_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_866_nl, CONVOLUTION_LOOP_for_for_for_for_mux_854_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_842_nl, CONVOLUTION_LOOP_for_for_for_for_mux_830_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_818_nl, CONVOLUTION_LOOP_for_for_for_for_mux_806_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_794_nl, CONVOLUTION_LOOP_for_for_for_for_mux_782_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_770_nl, CONVOLUTION_LOOP_for_for_for_for_mux_758_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_746_nl, CONVOLUTION_LOOP_for_for_for_for_mux_734_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_722_nl, CONVOLUTION_LOOP_for_for_for_for_mux_710_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_698_nl, CONVOLUTION_LOOP_for_for_for_for_mux_686_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_674_nl, CONVOLUTION_LOOP_for_for_for_for_mux_662_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_650_nl, CONVOLUTION_LOOP_for_for_for_for_mux_638_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_626_nl, CONVOLUTION_LOOP_for_for_for_for_mux_614_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_602_nl, CONVOLUTION_LOOP_for_for_for_for_mux_590_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_578_nl, CONVOLUTION_LOOP_for_for_for_for_mux_566_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_554_nl, CONVOLUTION_LOOP_for_for_for_for_mux_542_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_530_nl, CONVOLUTION_LOOP_for_for_for_for_mux_518_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_506_nl, CONVOLUTION_LOOP_for_for_for_for_mux_494_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_482_nl, CONVOLUTION_LOOP_for_for_for_for_mux_470_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_458_nl, CONVOLUTION_LOOP_for_for_for_for_mux_446_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_434_nl, CONVOLUTION_LOOP_for_for_for_for_mux_422_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_410_nl, CONVOLUTION_LOOP_for_for_for_for_mux_398_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_386_nl, CONVOLUTION_LOOP_for_for_for_for_mux_374_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_362_nl, CONVOLUTION_LOOP_for_for_for_for_mux_350_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_338_nl, CONVOLUTION_LOOP_for_for_for_for_mux_326_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_314_nl, CONVOLUTION_LOOP_for_for_for_for_mux_302_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_290_nl, CONVOLUTION_LOOP_for_for_for_for_mux_278_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_266_nl, CONVOLUTION_LOOP_for_for_for_for_mux_254_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_242_nl, CONVOLUTION_LOOP_for_for_for_for_mux_230_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_218_nl, CONVOLUTION_LOOP_for_for_for_for_mux_206_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_194_nl, CONVOLUTION_LOOP_for_for_for_for_mux_182_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_170_nl, CONVOLUTION_LOOP_for_for_for_for_mux_158_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_146_nl, CONVOLUTION_LOOP_for_for_for_for_mux_134_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_122_nl, CONVOLUTION_LOOP_for_for_for_for_mux_110_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_98_nl, CONVOLUTION_LOOP_for_for_for_for_mux_86_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_74_nl, CONVOLUTION_LOOP_for_for_for_for_mux_62_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_50_nl, CONVOLUTION_LOOP_for_for_for_for_mux_38_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_26_nl, CONVOLUTION_LOOP_for_for_for_for_mux_14_nl,
          CONVOLUTION_LOOP_for_for_for_for_mux_2_nl, {CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3
          , CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 , CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1_0});
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_2 <= CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1;
      CONVOLUTION_LOOP_for_for_for_unequal_tmp_1 <= (CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0!=5'b00000);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2
          <= 1'b0;
      exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_2 <= 1'b0;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_2 <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
          <= 1'b0;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
          <= 45'b000000000000000000000000000000000000000000000;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1
          <= 1'b0;
      exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      exit_COMPUTE_LOOP_lpi_1_dfm_2_st_2 <= 1'b0;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_if_1_and_6_cse ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_2
          <= CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1;
      exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_2 <= exit_CONVOLUTION_LOOP_lpi_1_dfm_3_st_1;
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_st_2 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_3_1;
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_itm_1
          <= CONVOLUTION_LOOP_for_for_for_acc_mux_5_nl & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_1_itm_1
          <= MUX_v_45_2_2(45'b000000000000000000000000000000000000000000000, CONVOLUTION_LOOP_for_for_for_acc_mux_3_nl,
          CONVOLUTION_LOOP_for_for_for_for_not_28_nl);
      CONVOLUTION_LOOP_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_and_2_itm_1
          <= CONVOLUTION_LOOP_for_for_for_acc_mux_1_nl & (~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1);
      exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_2 <= exitL_exit_CONVOLUTION_LOOP_lpi_1_dfm_st_1;
      exit_COMPUTE_LOOP_lpi_1_dfm_2_st_2 <= exit_COMPUTE_LOOP_lpi_1_dfm_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_3 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_2 <= 3'b000;
      n_w_out_lpi_1_dfm_1 <= 8'b00000000;
      n_h_out_lpi_1_dfm_1 <= 8'b00000000;
      COMPUTE_LOOP_b_4_0_lpi_1_3_0 <= 4'b0000;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 <= 3'b000;
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1_0 <= 1'b0;
      CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0 <= 5'b00000;
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1 <= 14'b00000000000000;
    end
    else if ( CONVOLUTION_LOOP_for_for_for_for_for_n_and_itm ) begin
      CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_3 <= MUX_v_3_2_2(CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_and_nl,
          CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_sva_2, or_277_nl);
      CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_2 <= MUX_v_3_2_2(CONVOLUTION_LOOP_for_for_for_for_m_2_0_sva_2,
          CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_4, and_74_nl);
      n_w_out_lpi_1_dfm_1 <= n_w_out_lpi_1_dfm_3;
      n_h_out_lpi_1_dfm_1 <= n_h_out_lpi_1_dfm_3;
      COMPUTE_LOOP_b_4_0_lpi_1_3_0 <= MUX_v_4_2_2((COMPUTE_LOOP_acc_tmp[3:0]), COMPUTE_LOOP_b_4_0_lpi_1_dfm_3_0_1,
          and_84_nl);
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3 <= nl_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3[4:0];
      CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_2_0 <= CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[2:0];
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_1_0 <= CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6[0];
      CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_1_4_0 <= CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0;
      CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1 <= nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1[13:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (and_131_cse | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_LOOP_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~(nand_tmp_7 | (~(or_113_cse & and_9_tmp)) | (fsm_output[0])))
        ) begin
      exit_COMPUTE_LOOP_sva_2 <= exit_COMPUTE_LOOP_sva_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_40 | or_dcpl_39 | (fsm_output[0]))) ) begin
      exit_CONVOLUTION_LOOP_lpi_1_dfm_1 <= or_113_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(mux_35_cse | or_dcpl_39 | (fsm_output[0]))) ) begin
      exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1 <= exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(mux_tmp_17 | not_tmp_22 | (~ and_9_tmp) | (fsm_output[0])))
        ) begin
      exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1 <= exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_66 | (~ and_9_tmp) | (fsm_output[0]))) ) begin
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1 <= exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_4_0 <= 5'b00000;
    end
    else if ( core_wen & (and_dcpl_72 | CONVOLUTION_LOOP_for_and_3_rgt | CONVOLUTION_LOOP_for_and_4_rgt)
        ) begin
      CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_4_0 <= MUX1HOT_v_5_3_2(({{4{or_113_cse}},
          or_113_cse}), (CONVOLUTION_LOOP_for_acc_tmp[4:0]), CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0,
          {and_dcpl_72 , CONVOLUTION_LOOP_for_and_3_rgt , CONVOLUTION_LOOP_for_and_4_rgt});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_2_4_0 <= 5'b00000;
    end
    else if ( core_wen & (and_dcpl_72 | and_dcpl_73) ) begin
      CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_2_4_0 <= MUX_v_5_2_2((CONVOLUTION_LOOP_acc_tmp[4:0]),
          CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_4_0_1, and_dcpl_73);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_4 <= 5'b00000;
    end
    else if ( core_wen & (and_88_rgt | CONVOLUTION_LOOP_for_for_and_3_rgt | CONVOLUTION_LOOP_for_for_and_4_rgt)
        ) begin
      CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_4 <= MUX1HOT_v_5_3_2(({{4{exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1_mx0w0}},
          exit_CONVOLUTION_LOOP_for_lpi_1_dfm_1_mx0w0}), CONVOLUTION_LOOP_for_for_i_4_0_sva_2,
          CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6, {and_88_rgt , CONVOLUTION_LOOP_for_for_and_3_rgt
          , CONVOLUTION_LOOP_for_for_and_4_rgt});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_4 <= 5'b00000;
    end
    else if ( core_wen & (and_90_rgt | CONVOLUTION_LOOP_for_for_for_and_2588_rgt
        | CONVOLUTION_LOOP_for_for_for_and_2589_rgt) ) begin
      CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_4 <= MUX1HOT_v_5_3_2(({{4{exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0}},
          exit_CONVOLUTION_LOOP_for_for_lpi_1_dfm_1_mx0w0}), CONVOLUTION_LOOP_for_for_for_j_4_0_sva_2,
          CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6, {and_90_rgt , CONVOLUTION_LOOP_for_for_for_and_2588_rgt
          , CONVOLUTION_LOOP_for_for_for_and_2589_rgt});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_1 <= 8'b00000000;
    end
    else if ( core_wen & (CONVOLUTION_LOOP_for_for_for_y_and_rgt | CONVOLUTION_LOOP_for_for_for_y_and_1_rgt
        | and_dcpl_59) ) begin
      CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_1 <= MUX1HOT_v_8_3_2(CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1,
          CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_1_dfm, z_out, {CONVOLUTION_LOOP_for_for_for_y_and_rgt
          , CONVOLUTION_LOOP_for_for_for_y_and_1_rgt , and_dcpl_59});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_1 <= 8'b00000000;
    end
    else if ( core_wen & (and_dcpl_57 | and_dcpl_59) ) begin
      CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_1 <= MUX_v_8_2_2(z_out, CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0,
          and_dcpl_59);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (((~ mux_tmp_17) & and_9_tmp & (fsm_output[1])) | CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1)
        ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1
          <= MUX_s_1_2_2(CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_if_CONVOLUTION_LOOP_for_if_nor_cse,
          CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm,
          CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm_1_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_1_dfm <= 8'b00000000;
    end
    else if ( core_wen & (~(and_dcpl_84 | (~ and_9_tmp))) ) begin
      CONVOLUTION_LOOP_for_for_for_y_mul_cse_lpi_1_dfm <= CONVOLUTION_LOOP_for_for_for_y_mul_cse_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm
          <= 1'b0;
    end
    else if ( core_wen & (~(mux_tmp_17 | (~ and_9_tmp) | (fsm_output[0]))) ) begin
      CONVOLUTION_LOOP_for_for_for_CONVOLUTION_LOOP_for_for_for_if_1_CONVOLUTION_LOOP_for_for_for_if_1_nor_itm
          <= CONVOLUTION_LOOP_for_CONVOLUTION_LOOP_for_if_CONVOLUTION_LOOP_for_if_nor_cse;
    end
  end
  assign or_89_nl = (operator_8_false_8_acc_tmp[8]) | COMPUTE_LOOP_if_COMPUTE_LOOP_if_nand_tmp
      | mux_tmp_21;
  assign mux_37_nl = MUX_s_1_2_2(or_89_nl, mux_tmp_21, COMPUTE_LOOP_acc_tmp[4]);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl = CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0
      * ({n_w_in_acc_psp_lpi_1_dfm_mx0 , conf_info_crt_lpi_1_dfm_192_mx0});
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_8_nl
      + conv_u2u_8_14(CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_mx0);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl = ({n_w_in_acc_psp_lpi_1_dfm_mx0
      , conf_info_crt_lpi_1_dfm_192_mx0}) * ({n_h_in_acc_psp_lpi_1_dfm_mx0 , conf_info_crt_lpi_1_dfm_160_mx0});
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_7_nl
      * CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0;
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_3_itm_1  = CONVOLUTION_LOOP_for_for_for_for_for_acc_12_nl
      + CONVOLUTION_LOOP_for_for_for_for_for_mul_6_nl;
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_4_nl = conv_u2u_13_13(CONVOLUTION_LOOP_for_k_5_0_lpi_1_dfm_4_0_mx0w0
      * conf_info_crt_lpi_1_dfm_103_96_mx0);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_4_nl
      * conf_info_crt_lpi_1_dfm_103_96_mx0;
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl[15:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_5_nl = conv_u2u_11_11(CONVOLUTION_LOOP_for_for_for_for_m_2_0_lpi_1_dfm_4
      * conf_info_crt_lpi_1_dfm_103_96_mx0);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_5_nl
      + conv_u2u_3_11(CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_5);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl[10:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_3_nl
      + conv_u2u_11_16(CONVOLUTION_LOOP_for_for_for_for_for_acc_10_nl);
  assign CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl[15:0];
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_2_nl = conv_u2u_13_13(CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_4_0_1
      * conf_info_crt_lpi_1_dfm_103_96_mx0);
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_1_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_2_nl
      * conf_info_crt_lpi_1_dfm_103_96_mx0;
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_1_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_1_nl[15:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_nl = CONVOLUTION_LOOP_for_for_for_for_for_mul_1_nl
      * conf_info_crt_lpi_1_dfm_135_128_mx0;
  assign CONVOLUTION_LOOP_for_for_for_for_for_mul_nl = nl_CONVOLUTION_LOOP_for_for_for_for_for_mul_nl[15:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_for_for_acc_itm_1  = CONVOLUTION_LOOP_for_for_for_for_for_acc_11_nl
      + CONVOLUTION_LOOP_for_for_for_for_for_mul_nl;
  assign CONVOLUTION_LOOP_for_for_for_for_mux_12_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_24_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_36_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_48_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_60_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_72_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_84_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_96_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_108_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_120_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_132_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_144_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_156_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_168_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_180_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_192_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_204_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_216_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_228_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_240_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_252_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_264_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_276_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_288_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_300_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_312_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_324_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_336_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_348_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_360_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_372_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_384_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_396_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_408_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_420_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_432_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_444_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_456_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_468_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_480_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_492_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_504_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_516_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_528_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_540_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_552_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_564_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_576_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_588_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_600_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_612_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_624_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_636_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_648_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_660_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_672_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_684_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_696_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_708_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_720_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_732_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_744_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_756_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_768_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_780_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_792_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_804_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_816_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_828_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_840_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_852_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_864_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_876_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_888_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_900_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_912_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_924_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_936_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_948_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_960_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_972_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_984_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_996_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1008_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1020_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1032_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1044_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1056_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1068_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1080_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1092_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1104_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1116_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1128_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1140_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1152_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1164_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1176_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1188_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1200_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1212_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1224_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1236_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1248_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1260_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1272_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1284_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1296_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1308_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1320_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1332_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1344_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1356_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1368_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1380_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1392_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1404_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1416_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1428_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1440_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1452_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1464_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1476_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1488_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1500_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1512_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1524_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1536_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1548_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1560_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1572_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1584_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1596_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1608_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1620_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1632_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1644_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1656_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1668_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1680_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1692_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1704_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1716_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1728_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1740_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1752_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1764_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1776_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1788_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1800_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1812_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1824_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1836_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1848_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1860_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1872_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1884_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1896_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1908_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1920_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1932_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1944_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1938_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1926_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1914_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1902_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1890_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1878_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1866_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1854_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1842_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1830_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1818_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1806_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1794_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1782_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1770_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1758_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1746_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1734_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1722_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1710_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1698_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1686_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1674_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1662_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1650_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1638_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1626_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1614_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1602_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1590_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1578_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1566_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1554_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1542_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1530_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1518_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1506_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1494_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1482_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1470_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1458_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1446_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1434_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1422_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1410_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1398_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1386_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1374_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1362_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1350_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1338_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1326_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1314_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1302_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1290_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1278_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1266_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1254_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1242_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1230_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1218_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1206_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1194_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1182_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1170_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1158_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1146_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1134_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1122_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1110_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1098_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1086_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1074_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1062_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1050_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1038_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1026_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1014_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1002_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_990_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_978_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_966_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_954_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_942_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_930_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_918_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_906_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_894_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_882_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_870_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_858_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_846_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_834_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_822_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_810_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_798_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_786_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_774_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_762_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_750_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_738_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_726_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_714_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_702_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_690_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_678_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_666_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_654_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_642_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_630_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_618_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_606_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_594_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_582_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_570_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_558_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_546_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_534_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_522_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_510_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_498_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_486_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_474_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_462_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_450_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_438_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_426_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_414_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_402_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_390_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_378_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_366_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_354_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_342_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_330_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_318_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_306_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_294_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_282_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_270_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_258_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_246_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_234_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_222_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_210_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_0_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_198_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_1_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_186_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_2_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_174_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_3_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_162_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_4_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_150_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_5_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_138_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_6_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_126_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_7_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_114_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_8_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_102_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_9_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_90_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_10_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_78_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_11_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_66_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_12_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_54_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_13_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_42_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_14_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_30_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_15_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_18_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_16_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_6_nl = MUX_v_11_2_2(COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_17_56_46_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_10_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_22_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_34_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_46_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_58_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_70_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_82_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_94_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_106_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_118_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_130_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_142_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_154_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_166_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_178_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_190_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_202_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_214_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_0_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_226_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_238_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_250_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_262_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_274_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_286_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_298_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_310_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_322_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_334_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_346_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_358_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_370_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_382_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_394_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_406_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_418_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_430_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_1_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_442_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_454_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_466_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_478_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_490_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_502_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_514_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_526_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_538_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_550_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_562_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_574_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_586_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_598_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_610_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_622_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_634_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_646_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_2_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_658_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_670_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_682_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_694_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_706_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_718_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_730_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_742_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_754_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_766_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_778_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_790_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_802_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_814_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_826_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_838_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_850_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_862_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_3_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_874_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_886_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_898_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_910_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_922_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_934_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_946_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_958_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_970_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_982_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_994_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1006_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1018_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1030_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1042_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1054_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1066_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1078_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_4_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1090_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1102_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1114_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1126_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1138_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1150_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1162_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1174_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1186_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1198_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1210_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1222_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1234_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1246_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1258_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1270_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1282_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1294_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_5_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1306_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1318_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1330_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1342_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1354_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1366_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1378_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1390_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1402_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1414_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1426_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1438_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1450_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1462_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1474_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1486_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1498_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1510_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_6_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1522_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1534_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1546_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1558_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1570_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1582_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1594_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1606_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1618_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1630_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1642_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1654_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1666_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1678_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1690_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1702_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1714_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1726_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_7_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1738_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1750_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1762_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1774_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1786_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1798_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1810_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1822_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1834_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1846_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1858_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1870_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1882_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1894_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1906_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1918_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1930_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1942_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_8_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1936_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1924_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1912_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1900_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1888_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1876_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1864_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1852_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1840_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1828_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1816_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1804_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1792_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1780_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1768_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1756_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1744_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1732_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_9_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1720_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1708_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1696_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1684_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1672_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1660_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1648_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1636_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1624_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1612_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1600_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1588_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1576_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1564_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1552_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1540_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1528_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1516_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_10_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1504_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1492_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1480_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1468_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1456_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1444_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1432_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1420_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1408_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1396_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1384_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1372_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1360_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1348_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1336_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1324_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1312_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1300_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_11_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1288_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1276_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1264_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1252_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1240_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1228_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1216_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1204_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1192_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1180_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1168_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1156_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1144_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1132_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1120_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1108_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1096_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1084_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_12_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1072_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1060_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1048_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1036_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1024_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1012_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1000_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_988_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_976_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_964_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_952_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_940_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_928_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_916_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_904_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_892_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_880_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_868_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_13_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_856_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_844_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_832_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_820_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_808_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_796_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_784_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_772_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_760_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_748_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_736_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_724_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_712_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_700_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_688_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_676_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_664_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_652_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_14_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_640_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_628_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_616_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_604_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_592_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_580_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_568_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_556_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_544_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_532_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_520_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_508_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_496_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_484_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_472_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_460_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_448_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_436_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_15_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_424_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_412_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_400_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_388_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_376_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_364_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_352_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_340_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_328_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_316_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_304_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_292_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_280_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_268_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_256_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_244_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_232_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_220_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_16_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_208_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_0_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_196_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_1_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_184_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_2_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_172_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_3_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_160_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_4_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_148_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_5_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_136_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_6_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_124_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_7_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_112_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_8_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_100_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_9_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_88_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_10_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_76_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_11_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_64_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_12_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_52_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_13_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_40_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_14_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_28_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_15_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_16_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_16_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_4_nl = MUX_v_45_2_2(COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_3,
      COMPUTE_LOOP_buf_acc_data_17_17_45_1_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_8_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_20_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_32_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_44_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_56_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_68_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_80_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_92_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_104_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_116_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_128_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_140_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_152_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_164_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_176_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_188_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_200_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_212_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_0_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_224_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_236_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_248_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_260_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_272_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_284_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_296_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_308_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_320_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_332_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_344_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_356_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_368_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_380_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_392_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_404_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_416_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_428_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_1_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_440_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_452_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_464_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_476_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_488_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_500_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_512_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_524_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_536_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_548_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_560_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_572_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_584_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_596_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_608_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_620_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_632_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_644_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_2_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_656_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_668_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_680_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_692_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_704_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_716_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_728_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_740_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_752_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_764_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_776_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_788_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_800_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_812_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_824_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_836_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_848_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_860_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_3_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_872_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_884_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_896_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_908_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_920_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_932_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_944_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_956_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_968_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_980_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_992_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1004_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1016_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1028_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1040_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1052_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1064_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1076_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_4_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1088_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1100_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1112_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1124_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1136_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1148_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1160_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1172_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1184_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1196_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1208_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1220_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1232_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1244_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1256_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1268_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1280_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1292_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_5_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1304_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1316_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1328_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1340_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1352_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1364_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1376_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1388_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1400_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1412_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1424_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1436_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1448_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1460_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1472_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1484_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1496_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1508_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_6_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1520_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1532_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1544_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1556_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1568_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1580_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1592_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1604_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1616_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1628_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1640_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1652_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1664_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1676_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1688_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1700_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1712_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1724_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_7_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1736_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1748_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1760_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1772_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1784_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1796_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1808_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1820_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1832_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1844_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1856_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1868_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1880_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1892_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1904_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1916_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1928_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1940_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_8_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1934_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1922_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1910_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1898_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1886_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1874_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1862_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1850_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1838_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1826_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1814_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1802_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1790_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1778_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1766_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1754_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1742_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1730_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_9_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1718_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1706_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1694_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1682_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1670_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1658_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1646_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1634_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1622_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1610_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1598_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1586_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1574_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1562_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1550_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1538_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1526_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1514_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_10_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1502_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1490_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1478_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1466_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1454_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1442_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1430_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1418_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1406_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1394_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1382_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1370_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1358_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1346_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1334_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1322_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1310_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1298_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_11_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1286_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1274_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1262_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1250_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1238_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1226_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1214_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1202_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1190_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1178_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1166_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1154_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1142_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1130_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1118_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1106_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1094_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1082_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_12_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1070_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1058_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1046_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1034_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1022_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_1010_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_998_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_986_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_974_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_962_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_950_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_938_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_926_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_914_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_902_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_890_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_878_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_866_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_13_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_854_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_842_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_830_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_818_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_806_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_794_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_782_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_770_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_758_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_746_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_734_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_722_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_710_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_698_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_686_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_674_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_662_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_650_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_14_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_638_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_626_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_614_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_602_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_590_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_578_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_566_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_554_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_542_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_530_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_518_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_506_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_494_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_482_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_470_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_458_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_446_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_434_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_15_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_422_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_410_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_398_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_386_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_374_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_362_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_350_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_338_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_326_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_314_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_302_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_290_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_278_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_266_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_254_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_242_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_230_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_218_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_16_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_206_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_0_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_194_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_1_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_182_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_2_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_170_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_3_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_158_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_4_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_146_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_5_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_134_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_6_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_122_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_7_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_110_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_8_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_98_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_9_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_86_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_10_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_74_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_11_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_62_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_12_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_50_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_13_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_38_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_14_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_26_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_15_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_14_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_16_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_for_mux_2_nl = MUX_s_1_2_2(COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_1_mx0,
      COMPUTE_LOOP_buf_acc_data_17_17_0_lpi_1_dfm_2, or_dcpl_31);
  assign CONVOLUTION_LOOP_for_for_for_acc_mux_5_nl = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_46_sva_1,
      CONVOLUTION_LOOP_for_for_for_acc_46_sva_1_mx0w0, and_5_tmp);
  assign CONVOLUTION_LOOP_for_for_for_acc_mux_3_nl = MUX_v_45_2_2(CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1,
      CONVOLUTION_LOOP_for_for_for_acc_45_1_sva_1_mx0w0, and_5_tmp);
  assign CONVOLUTION_LOOP_for_for_for_for_not_28_nl = ~ exitL_exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1;
  assign CONVOLUTION_LOOP_for_for_for_acc_mux_1_nl = MUX_s_1_2_2(CONVOLUTION_LOOP_for_for_for_acc_0_sva_1,
      CONVOLUTION_LOOP_for_for_for_acc_0_sva_1_mx0w0, and_5_tmp);
  assign CONVOLUTION_LOOP_for_for_for_for_for_CONVOLUTION_LOOP_for_for_for_for_for_and_nl
      = MUX_v_3_2_2(3'b000, CONVOLUTION_LOOP_for_for_for_for_for_n_2_0_lpi_1_dfm_5,
      exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0);
  assign or_277_nl = (and_dcpl_57 & exit_CONVOLUTION_LOOP_for_for_for_for_lpi_1_dfm_1_mx0w0
      & or_dcpl_34) | and_dcpl_59;
  assign nor_51_nl = ~((~ CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp) | CONVOLUTION_LOOP_for_for_for_for_if_equal_tmp
      | (~ CONVOLUTION_LOOP_for_for_for_for_for_if_nor_tmp) | (operator_8_false_1_acc_tmp[8]));
  assign mux_65_nl = MUX_s_1_2_2(or_73_cse, nor_51_nl, operator_8_false_6_acc_itm_3_1);
  assign and_74_nl = (~ mux_65_nl) & and_9_tmp;
  assign and_84_nl = mux_tmp_21 & and_9_tmp;
  assign nl_CONVOLUTION_LOOP_for_for_for_else_acc_psp_sva_1_7_3  = conv_u2u_2_5(CONVOLUTION_LOOP_for_for_for_if_acc_1_ncse_1[4:3])
      + CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6;
  assign CONVOLUTION_LOOP_for_for_for_index_out_mul_2_nl = conv_u2u_13_13(CONVOLUTION_LOOP_for_for_i_4_0_lpi_1_dfm_6
      * n_w_out_lpi_1_dfm_3);
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl = CONVOLUTION_LOOP_for_for_for_index_out_mul_2_nl
      + conv_u2u_5_13(CONVOLUTION_LOOP_for_for_for_j_4_0_lpi_1_dfm_6);
  assign CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl = nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl[12:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl = n_w_out_lpi_1_dfm_3
      * n_h_out_lpi_1_dfm_3;
  assign CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl = nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_nl = CONVOLUTION_LOOP_for_for_for_index_out_mul_1_nl
      * CONVOLUTION_LOOP_fl_5_0_lpi_1_dfm_4_0_1;
  assign CONVOLUTION_LOOP_for_for_for_index_out_mul_nl = nl_CONVOLUTION_LOOP_for_for_for_index_out_mul_nl[13:0];
  assign nl_CONVOLUTION_LOOP_for_for_for_index_out_acc_itm_1  = conv_u2u_13_14(CONVOLUTION_LOOP_for_for_for_index_out_acc_2_nl)
      + CONVOLUTION_LOOP_for_for_for_index_out_mul_nl;
  assign and_275_nl = (~((~((operator_8_false_1_acc_tmp[8:3]==6'b000000) & CONVOLUTION_LOOP_for_for_for_for_for_if_equal_tmp))
      & operator_8_false_6_acc_itm_3_1)) & (fsm_output[1]);
  assign CONVOLUTION_LOOP_for_for_for_for_for_mux_6_nl = MUX_v_8_2_2(CONVOLUTION_LOOP_for_for_for_y_lpi_1_dfm_mx0,
      CONVOLUTION_LOOP_for_for_for_x_lpi_1_dfm_mx0, and_275_nl);
  assign nl_z_out = CONVOLUTION_LOOP_for_for_for_for_for_mux_6_nl + 8'b00000001;
  assign z_out = nl_z_out[7:0];

  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [44:0] MUX1HOT_v_45_3_2;
    input [44:0] input_2;
    input [44:0] input_1;
    input [44:0] input_0;
    input [2:0] sel;
    reg [44:0] result;
  begin
    result = input_0 & {45{sel[0]}};
    result = result | ( input_1 & {45{sel[1]}});
    result = result | ( input_2 & {45{sel[2]}});
    MUX1HOT_v_45_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_324_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] input_2;
    input [0:0] input_3;
    input [0:0] input_4;
    input [0:0] input_5;
    input [0:0] input_6;
    input [0:0] input_7;
    input [0:0] input_8;
    input [0:0] input_9;
    input [0:0] input_10;
    input [0:0] input_11;
    input [0:0] input_12;
    input [0:0] input_13;
    input [0:0] input_14;
    input [0:0] input_15;
    input [0:0] input_16;
    input [0:0] input_17;
    input [0:0] input_18;
    input [0:0] input_19;
    input [0:0] input_20;
    input [0:0] input_21;
    input [0:0] input_22;
    input [0:0] input_23;
    input [0:0] input_24;
    input [0:0] input_25;
    input [0:0] input_26;
    input [0:0] input_27;
    input [0:0] input_28;
    input [0:0] input_29;
    input [0:0] input_30;
    input [0:0] input_31;
    input [0:0] input_32;
    input [0:0] input_33;
    input [0:0] input_34;
    input [0:0] input_35;
    input [0:0] input_36;
    input [0:0] input_37;
    input [0:0] input_38;
    input [0:0] input_39;
    input [0:0] input_40;
    input [0:0] input_41;
    input [0:0] input_42;
    input [0:0] input_43;
    input [0:0] input_44;
    input [0:0] input_45;
    input [0:0] input_46;
    input [0:0] input_47;
    input [0:0] input_48;
    input [0:0] input_49;
    input [0:0] input_50;
    input [0:0] input_51;
    input [0:0] input_52;
    input [0:0] input_53;
    input [0:0] input_54;
    input [0:0] input_55;
    input [0:0] input_56;
    input [0:0] input_57;
    input [0:0] input_58;
    input [0:0] input_59;
    input [0:0] input_60;
    input [0:0] input_61;
    input [0:0] input_62;
    input [0:0] input_63;
    input [0:0] input_64;
    input [0:0] input_65;
    input [0:0] input_66;
    input [0:0] input_67;
    input [0:0] input_68;
    input [0:0] input_69;
    input [0:0] input_70;
    input [0:0] input_71;
    input [0:0] input_72;
    input [0:0] input_73;
    input [0:0] input_74;
    input [0:0] input_75;
    input [0:0] input_76;
    input [0:0] input_77;
    input [0:0] input_78;
    input [0:0] input_79;
    input [0:0] input_80;
    input [0:0] input_81;
    input [0:0] input_82;
    input [0:0] input_83;
    input [0:0] input_84;
    input [0:0] input_85;
    input [0:0] input_86;
    input [0:0] input_87;
    input [0:0] input_88;
    input [0:0] input_89;
    input [0:0] input_90;
    input [0:0] input_91;
    input [0:0] input_92;
    input [0:0] input_93;
    input [0:0] input_94;
    input [0:0] input_95;
    input [0:0] input_96;
    input [0:0] input_97;
    input [0:0] input_98;
    input [0:0] input_99;
    input [0:0] input_100;
    input [0:0] input_101;
    input [0:0] input_102;
    input [0:0] input_103;
    input [0:0] input_104;
    input [0:0] input_105;
    input [0:0] input_106;
    input [0:0] input_107;
    input [0:0] input_108;
    input [0:0] input_109;
    input [0:0] input_110;
    input [0:0] input_111;
    input [0:0] input_112;
    input [0:0] input_113;
    input [0:0] input_114;
    input [0:0] input_115;
    input [0:0] input_116;
    input [0:0] input_117;
    input [0:0] input_118;
    input [0:0] input_119;
    input [0:0] input_120;
    input [0:0] input_121;
    input [0:0] input_122;
    input [0:0] input_123;
    input [0:0] input_124;
    input [0:0] input_125;
    input [0:0] input_126;
    input [0:0] input_127;
    input [0:0] input_128;
    input [0:0] input_129;
    input [0:0] input_130;
    input [0:0] input_131;
    input [0:0] input_132;
    input [0:0] input_133;
    input [0:0] input_134;
    input [0:0] input_135;
    input [0:0] input_136;
    input [0:0] input_137;
    input [0:0] input_138;
    input [0:0] input_139;
    input [0:0] input_140;
    input [0:0] input_141;
    input [0:0] input_142;
    input [0:0] input_143;
    input [0:0] input_144;
    input [0:0] input_145;
    input [0:0] input_146;
    input [0:0] input_147;
    input [0:0] input_148;
    input [0:0] input_149;
    input [0:0] input_150;
    input [0:0] input_151;
    input [0:0] input_152;
    input [0:0] input_153;
    input [0:0] input_154;
    input [0:0] input_155;
    input [0:0] input_156;
    input [0:0] input_157;
    input [0:0] input_158;
    input [0:0] input_159;
    input [0:0] input_160;
    input [0:0] input_161;
    input [0:0] input_162;
    input [0:0] input_163;
    input [0:0] input_164;
    input [0:0] input_165;
    input [0:0] input_166;
    input [0:0] input_167;
    input [0:0] input_168;
    input [0:0] input_169;
    input [0:0] input_170;
    input [0:0] input_171;
    input [0:0] input_172;
    input [0:0] input_173;
    input [0:0] input_174;
    input [0:0] input_175;
    input [0:0] input_176;
    input [0:0] input_177;
    input [0:0] input_178;
    input [0:0] input_179;
    input [0:0] input_180;
    input [0:0] input_181;
    input [0:0] input_182;
    input [0:0] input_183;
    input [0:0] input_184;
    input [0:0] input_185;
    input [0:0] input_186;
    input [0:0] input_187;
    input [0:0] input_188;
    input [0:0] input_189;
    input [0:0] input_190;
    input [0:0] input_191;
    input [0:0] input_192;
    input [0:0] input_193;
    input [0:0] input_194;
    input [0:0] input_195;
    input [0:0] input_196;
    input [0:0] input_197;
    input [0:0] input_198;
    input [0:0] input_199;
    input [0:0] input_200;
    input [0:0] input_201;
    input [0:0] input_202;
    input [0:0] input_203;
    input [0:0] input_204;
    input [0:0] input_205;
    input [0:0] input_206;
    input [0:0] input_207;
    input [0:0] input_208;
    input [0:0] input_209;
    input [0:0] input_210;
    input [0:0] input_211;
    input [0:0] input_212;
    input [0:0] input_213;
    input [0:0] input_214;
    input [0:0] input_215;
    input [0:0] input_216;
    input [0:0] input_217;
    input [0:0] input_218;
    input [0:0] input_219;
    input [0:0] input_220;
    input [0:0] input_221;
    input [0:0] input_222;
    input [0:0] input_223;
    input [0:0] input_224;
    input [0:0] input_225;
    input [0:0] input_226;
    input [0:0] input_227;
    input [0:0] input_228;
    input [0:0] input_229;
    input [0:0] input_230;
    input [0:0] input_231;
    input [0:0] input_232;
    input [0:0] input_233;
    input [0:0] input_234;
    input [0:0] input_235;
    input [0:0] input_236;
    input [0:0] input_237;
    input [0:0] input_238;
    input [0:0] input_239;
    input [0:0] input_240;
    input [0:0] input_241;
    input [0:0] input_242;
    input [0:0] input_243;
    input [0:0] input_244;
    input [0:0] input_245;
    input [0:0] input_246;
    input [0:0] input_247;
    input [0:0] input_248;
    input [0:0] input_249;
    input [0:0] input_250;
    input [0:0] input_251;
    input [0:0] input_252;
    input [0:0] input_253;
    input [0:0] input_254;
    input [0:0] input_255;
    input [0:0] input_256;
    input [0:0] input_257;
    input [0:0] input_258;
    input [0:0] input_259;
    input [0:0] input_260;
    input [0:0] input_261;
    input [0:0] input_262;
    input [0:0] input_263;
    input [0:0] input_264;
    input [0:0] input_265;
    input [0:0] input_266;
    input [0:0] input_267;
    input [0:0] input_268;
    input [0:0] input_269;
    input [0:0] input_270;
    input [0:0] input_271;
    input [0:0] input_272;
    input [0:0] input_273;
    input [0:0] input_274;
    input [0:0] input_275;
    input [0:0] input_276;
    input [0:0] input_277;
    input [0:0] input_278;
    input [0:0] input_279;
    input [0:0] input_280;
    input [0:0] input_281;
    input [0:0] input_282;
    input [0:0] input_283;
    input [0:0] input_284;
    input [0:0] input_285;
    input [0:0] input_286;
    input [0:0] input_287;
    input [0:0] input_288;
    input [0:0] input_289;
    input [0:0] input_290;
    input [0:0] input_291;
    input [0:0] input_292;
    input [0:0] input_293;
    input [0:0] input_294;
    input [0:0] input_295;
    input [0:0] input_296;
    input [0:0] input_297;
    input [0:0] input_298;
    input [0:0] input_299;
    input [0:0] input_300;
    input [0:0] input_301;
    input [0:0] input_302;
    input [0:0] input_303;
    input [0:0] input_304;
    input [0:0] input_305;
    input [0:0] input_306;
    input [0:0] input_307;
    input [0:0] input_308;
    input [0:0] input_309;
    input [0:0] input_310;
    input [0:0] input_311;
    input [0:0] input_312;
    input [0:0] input_313;
    input [0:0] input_314;
    input [0:0] input_315;
    input [0:0] input_316;
    input [0:0] input_317;
    input [0:0] input_318;
    input [0:0] input_319;
    input [0:0] input_320;
    input [0:0] input_321;
    input [0:0] input_322;
    input [0:0] input_323;
    input [8:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_s_1_324_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_324_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [10:0] input_8;
    input [10:0] input_9;
    input [10:0] input_10;
    input [10:0] input_11;
    input [10:0] input_12;
    input [10:0] input_13;
    input [10:0] input_14;
    input [10:0] input_15;
    input [10:0] input_16;
    input [10:0] input_17;
    input [10:0] input_18;
    input [10:0] input_19;
    input [10:0] input_20;
    input [10:0] input_21;
    input [10:0] input_22;
    input [10:0] input_23;
    input [10:0] input_24;
    input [10:0] input_25;
    input [10:0] input_26;
    input [10:0] input_27;
    input [10:0] input_28;
    input [10:0] input_29;
    input [10:0] input_30;
    input [10:0] input_31;
    input [10:0] input_32;
    input [10:0] input_33;
    input [10:0] input_34;
    input [10:0] input_35;
    input [10:0] input_36;
    input [10:0] input_37;
    input [10:0] input_38;
    input [10:0] input_39;
    input [10:0] input_40;
    input [10:0] input_41;
    input [10:0] input_42;
    input [10:0] input_43;
    input [10:0] input_44;
    input [10:0] input_45;
    input [10:0] input_46;
    input [10:0] input_47;
    input [10:0] input_48;
    input [10:0] input_49;
    input [10:0] input_50;
    input [10:0] input_51;
    input [10:0] input_52;
    input [10:0] input_53;
    input [10:0] input_54;
    input [10:0] input_55;
    input [10:0] input_56;
    input [10:0] input_57;
    input [10:0] input_58;
    input [10:0] input_59;
    input [10:0] input_60;
    input [10:0] input_61;
    input [10:0] input_62;
    input [10:0] input_63;
    input [10:0] input_64;
    input [10:0] input_65;
    input [10:0] input_66;
    input [10:0] input_67;
    input [10:0] input_68;
    input [10:0] input_69;
    input [10:0] input_70;
    input [10:0] input_71;
    input [10:0] input_72;
    input [10:0] input_73;
    input [10:0] input_74;
    input [10:0] input_75;
    input [10:0] input_76;
    input [10:0] input_77;
    input [10:0] input_78;
    input [10:0] input_79;
    input [10:0] input_80;
    input [10:0] input_81;
    input [10:0] input_82;
    input [10:0] input_83;
    input [10:0] input_84;
    input [10:0] input_85;
    input [10:0] input_86;
    input [10:0] input_87;
    input [10:0] input_88;
    input [10:0] input_89;
    input [10:0] input_90;
    input [10:0] input_91;
    input [10:0] input_92;
    input [10:0] input_93;
    input [10:0] input_94;
    input [10:0] input_95;
    input [10:0] input_96;
    input [10:0] input_97;
    input [10:0] input_98;
    input [10:0] input_99;
    input [10:0] input_100;
    input [10:0] input_101;
    input [10:0] input_102;
    input [10:0] input_103;
    input [10:0] input_104;
    input [10:0] input_105;
    input [10:0] input_106;
    input [10:0] input_107;
    input [10:0] input_108;
    input [10:0] input_109;
    input [10:0] input_110;
    input [10:0] input_111;
    input [10:0] input_112;
    input [10:0] input_113;
    input [10:0] input_114;
    input [10:0] input_115;
    input [10:0] input_116;
    input [10:0] input_117;
    input [10:0] input_118;
    input [10:0] input_119;
    input [10:0] input_120;
    input [10:0] input_121;
    input [10:0] input_122;
    input [10:0] input_123;
    input [10:0] input_124;
    input [10:0] input_125;
    input [10:0] input_126;
    input [10:0] input_127;
    input [10:0] input_128;
    input [10:0] input_129;
    input [10:0] input_130;
    input [10:0] input_131;
    input [10:0] input_132;
    input [10:0] input_133;
    input [10:0] input_134;
    input [10:0] input_135;
    input [10:0] input_136;
    input [10:0] input_137;
    input [10:0] input_138;
    input [10:0] input_139;
    input [10:0] input_140;
    input [10:0] input_141;
    input [10:0] input_142;
    input [10:0] input_143;
    input [10:0] input_144;
    input [10:0] input_145;
    input [10:0] input_146;
    input [10:0] input_147;
    input [10:0] input_148;
    input [10:0] input_149;
    input [10:0] input_150;
    input [10:0] input_151;
    input [10:0] input_152;
    input [10:0] input_153;
    input [10:0] input_154;
    input [10:0] input_155;
    input [10:0] input_156;
    input [10:0] input_157;
    input [10:0] input_158;
    input [10:0] input_159;
    input [10:0] input_160;
    input [10:0] input_161;
    input [10:0] input_162;
    input [10:0] input_163;
    input [10:0] input_164;
    input [10:0] input_165;
    input [10:0] input_166;
    input [10:0] input_167;
    input [10:0] input_168;
    input [10:0] input_169;
    input [10:0] input_170;
    input [10:0] input_171;
    input [10:0] input_172;
    input [10:0] input_173;
    input [10:0] input_174;
    input [10:0] input_175;
    input [10:0] input_176;
    input [10:0] input_177;
    input [10:0] input_178;
    input [10:0] input_179;
    input [10:0] input_180;
    input [10:0] input_181;
    input [10:0] input_182;
    input [10:0] input_183;
    input [10:0] input_184;
    input [10:0] input_185;
    input [10:0] input_186;
    input [10:0] input_187;
    input [10:0] input_188;
    input [10:0] input_189;
    input [10:0] input_190;
    input [10:0] input_191;
    input [10:0] input_192;
    input [10:0] input_193;
    input [10:0] input_194;
    input [10:0] input_195;
    input [10:0] input_196;
    input [10:0] input_197;
    input [10:0] input_198;
    input [10:0] input_199;
    input [10:0] input_200;
    input [10:0] input_201;
    input [10:0] input_202;
    input [10:0] input_203;
    input [10:0] input_204;
    input [10:0] input_205;
    input [10:0] input_206;
    input [10:0] input_207;
    input [10:0] input_208;
    input [10:0] input_209;
    input [10:0] input_210;
    input [10:0] input_211;
    input [10:0] input_212;
    input [10:0] input_213;
    input [10:0] input_214;
    input [10:0] input_215;
    input [10:0] input_216;
    input [10:0] input_217;
    input [10:0] input_218;
    input [10:0] input_219;
    input [10:0] input_220;
    input [10:0] input_221;
    input [10:0] input_222;
    input [10:0] input_223;
    input [10:0] input_224;
    input [10:0] input_225;
    input [10:0] input_226;
    input [10:0] input_227;
    input [10:0] input_228;
    input [10:0] input_229;
    input [10:0] input_230;
    input [10:0] input_231;
    input [10:0] input_232;
    input [10:0] input_233;
    input [10:0] input_234;
    input [10:0] input_235;
    input [10:0] input_236;
    input [10:0] input_237;
    input [10:0] input_238;
    input [10:0] input_239;
    input [10:0] input_240;
    input [10:0] input_241;
    input [10:0] input_242;
    input [10:0] input_243;
    input [10:0] input_244;
    input [10:0] input_245;
    input [10:0] input_246;
    input [10:0] input_247;
    input [10:0] input_248;
    input [10:0] input_249;
    input [10:0] input_250;
    input [10:0] input_251;
    input [10:0] input_252;
    input [10:0] input_253;
    input [10:0] input_254;
    input [10:0] input_255;
    input [10:0] input_256;
    input [10:0] input_257;
    input [10:0] input_258;
    input [10:0] input_259;
    input [10:0] input_260;
    input [10:0] input_261;
    input [10:0] input_262;
    input [10:0] input_263;
    input [10:0] input_264;
    input [10:0] input_265;
    input [10:0] input_266;
    input [10:0] input_267;
    input [10:0] input_268;
    input [10:0] input_269;
    input [10:0] input_270;
    input [10:0] input_271;
    input [10:0] input_272;
    input [10:0] input_273;
    input [10:0] input_274;
    input [10:0] input_275;
    input [10:0] input_276;
    input [10:0] input_277;
    input [10:0] input_278;
    input [10:0] input_279;
    input [10:0] input_280;
    input [10:0] input_281;
    input [10:0] input_282;
    input [10:0] input_283;
    input [10:0] input_284;
    input [10:0] input_285;
    input [10:0] input_286;
    input [10:0] input_287;
    input [10:0] input_288;
    input [10:0] input_289;
    input [10:0] input_290;
    input [10:0] input_291;
    input [10:0] input_292;
    input [10:0] input_293;
    input [10:0] input_294;
    input [10:0] input_295;
    input [10:0] input_296;
    input [10:0] input_297;
    input [10:0] input_298;
    input [10:0] input_299;
    input [10:0] input_300;
    input [10:0] input_301;
    input [10:0] input_302;
    input [10:0] input_303;
    input [10:0] input_304;
    input [10:0] input_305;
    input [10:0] input_306;
    input [10:0] input_307;
    input [10:0] input_308;
    input [10:0] input_309;
    input [10:0] input_310;
    input [10:0] input_311;
    input [10:0] input_312;
    input [10:0] input_313;
    input [10:0] input_314;
    input [10:0] input_315;
    input [10:0] input_316;
    input [10:0] input_317;
    input [10:0] input_318;
    input [10:0] input_319;
    input [10:0] input_320;
    input [10:0] input_321;
    input [10:0] input_322;
    input [10:0] input_323;
    input [8:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_v_11_324_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [44:0] MUX_v_45_2_2;
    input [44:0] input_0;
    input [44:0] input_1;
    input [0:0] sel;
    reg [44:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_45_2_2 = result;
  end
  endfunction


  function automatic [44:0] MUX_v_45_324_2;
    input [44:0] input_0;
    input [44:0] input_1;
    input [44:0] input_2;
    input [44:0] input_3;
    input [44:0] input_4;
    input [44:0] input_5;
    input [44:0] input_6;
    input [44:0] input_7;
    input [44:0] input_8;
    input [44:0] input_9;
    input [44:0] input_10;
    input [44:0] input_11;
    input [44:0] input_12;
    input [44:0] input_13;
    input [44:0] input_14;
    input [44:0] input_15;
    input [44:0] input_16;
    input [44:0] input_17;
    input [44:0] input_18;
    input [44:0] input_19;
    input [44:0] input_20;
    input [44:0] input_21;
    input [44:0] input_22;
    input [44:0] input_23;
    input [44:0] input_24;
    input [44:0] input_25;
    input [44:0] input_26;
    input [44:0] input_27;
    input [44:0] input_28;
    input [44:0] input_29;
    input [44:0] input_30;
    input [44:0] input_31;
    input [44:0] input_32;
    input [44:0] input_33;
    input [44:0] input_34;
    input [44:0] input_35;
    input [44:0] input_36;
    input [44:0] input_37;
    input [44:0] input_38;
    input [44:0] input_39;
    input [44:0] input_40;
    input [44:0] input_41;
    input [44:0] input_42;
    input [44:0] input_43;
    input [44:0] input_44;
    input [44:0] input_45;
    input [44:0] input_46;
    input [44:0] input_47;
    input [44:0] input_48;
    input [44:0] input_49;
    input [44:0] input_50;
    input [44:0] input_51;
    input [44:0] input_52;
    input [44:0] input_53;
    input [44:0] input_54;
    input [44:0] input_55;
    input [44:0] input_56;
    input [44:0] input_57;
    input [44:0] input_58;
    input [44:0] input_59;
    input [44:0] input_60;
    input [44:0] input_61;
    input [44:0] input_62;
    input [44:0] input_63;
    input [44:0] input_64;
    input [44:0] input_65;
    input [44:0] input_66;
    input [44:0] input_67;
    input [44:0] input_68;
    input [44:0] input_69;
    input [44:0] input_70;
    input [44:0] input_71;
    input [44:0] input_72;
    input [44:0] input_73;
    input [44:0] input_74;
    input [44:0] input_75;
    input [44:0] input_76;
    input [44:0] input_77;
    input [44:0] input_78;
    input [44:0] input_79;
    input [44:0] input_80;
    input [44:0] input_81;
    input [44:0] input_82;
    input [44:0] input_83;
    input [44:0] input_84;
    input [44:0] input_85;
    input [44:0] input_86;
    input [44:0] input_87;
    input [44:0] input_88;
    input [44:0] input_89;
    input [44:0] input_90;
    input [44:0] input_91;
    input [44:0] input_92;
    input [44:0] input_93;
    input [44:0] input_94;
    input [44:0] input_95;
    input [44:0] input_96;
    input [44:0] input_97;
    input [44:0] input_98;
    input [44:0] input_99;
    input [44:0] input_100;
    input [44:0] input_101;
    input [44:0] input_102;
    input [44:0] input_103;
    input [44:0] input_104;
    input [44:0] input_105;
    input [44:0] input_106;
    input [44:0] input_107;
    input [44:0] input_108;
    input [44:0] input_109;
    input [44:0] input_110;
    input [44:0] input_111;
    input [44:0] input_112;
    input [44:0] input_113;
    input [44:0] input_114;
    input [44:0] input_115;
    input [44:0] input_116;
    input [44:0] input_117;
    input [44:0] input_118;
    input [44:0] input_119;
    input [44:0] input_120;
    input [44:0] input_121;
    input [44:0] input_122;
    input [44:0] input_123;
    input [44:0] input_124;
    input [44:0] input_125;
    input [44:0] input_126;
    input [44:0] input_127;
    input [44:0] input_128;
    input [44:0] input_129;
    input [44:0] input_130;
    input [44:0] input_131;
    input [44:0] input_132;
    input [44:0] input_133;
    input [44:0] input_134;
    input [44:0] input_135;
    input [44:0] input_136;
    input [44:0] input_137;
    input [44:0] input_138;
    input [44:0] input_139;
    input [44:0] input_140;
    input [44:0] input_141;
    input [44:0] input_142;
    input [44:0] input_143;
    input [44:0] input_144;
    input [44:0] input_145;
    input [44:0] input_146;
    input [44:0] input_147;
    input [44:0] input_148;
    input [44:0] input_149;
    input [44:0] input_150;
    input [44:0] input_151;
    input [44:0] input_152;
    input [44:0] input_153;
    input [44:0] input_154;
    input [44:0] input_155;
    input [44:0] input_156;
    input [44:0] input_157;
    input [44:0] input_158;
    input [44:0] input_159;
    input [44:0] input_160;
    input [44:0] input_161;
    input [44:0] input_162;
    input [44:0] input_163;
    input [44:0] input_164;
    input [44:0] input_165;
    input [44:0] input_166;
    input [44:0] input_167;
    input [44:0] input_168;
    input [44:0] input_169;
    input [44:0] input_170;
    input [44:0] input_171;
    input [44:0] input_172;
    input [44:0] input_173;
    input [44:0] input_174;
    input [44:0] input_175;
    input [44:0] input_176;
    input [44:0] input_177;
    input [44:0] input_178;
    input [44:0] input_179;
    input [44:0] input_180;
    input [44:0] input_181;
    input [44:0] input_182;
    input [44:0] input_183;
    input [44:0] input_184;
    input [44:0] input_185;
    input [44:0] input_186;
    input [44:0] input_187;
    input [44:0] input_188;
    input [44:0] input_189;
    input [44:0] input_190;
    input [44:0] input_191;
    input [44:0] input_192;
    input [44:0] input_193;
    input [44:0] input_194;
    input [44:0] input_195;
    input [44:0] input_196;
    input [44:0] input_197;
    input [44:0] input_198;
    input [44:0] input_199;
    input [44:0] input_200;
    input [44:0] input_201;
    input [44:0] input_202;
    input [44:0] input_203;
    input [44:0] input_204;
    input [44:0] input_205;
    input [44:0] input_206;
    input [44:0] input_207;
    input [44:0] input_208;
    input [44:0] input_209;
    input [44:0] input_210;
    input [44:0] input_211;
    input [44:0] input_212;
    input [44:0] input_213;
    input [44:0] input_214;
    input [44:0] input_215;
    input [44:0] input_216;
    input [44:0] input_217;
    input [44:0] input_218;
    input [44:0] input_219;
    input [44:0] input_220;
    input [44:0] input_221;
    input [44:0] input_222;
    input [44:0] input_223;
    input [44:0] input_224;
    input [44:0] input_225;
    input [44:0] input_226;
    input [44:0] input_227;
    input [44:0] input_228;
    input [44:0] input_229;
    input [44:0] input_230;
    input [44:0] input_231;
    input [44:0] input_232;
    input [44:0] input_233;
    input [44:0] input_234;
    input [44:0] input_235;
    input [44:0] input_236;
    input [44:0] input_237;
    input [44:0] input_238;
    input [44:0] input_239;
    input [44:0] input_240;
    input [44:0] input_241;
    input [44:0] input_242;
    input [44:0] input_243;
    input [44:0] input_244;
    input [44:0] input_245;
    input [44:0] input_246;
    input [44:0] input_247;
    input [44:0] input_248;
    input [44:0] input_249;
    input [44:0] input_250;
    input [44:0] input_251;
    input [44:0] input_252;
    input [44:0] input_253;
    input [44:0] input_254;
    input [44:0] input_255;
    input [44:0] input_256;
    input [44:0] input_257;
    input [44:0] input_258;
    input [44:0] input_259;
    input [44:0] input_260;
    input [44:0] input_261;
    input [44:0] input_262;
    input [44:0] input_263;
    input [44:0] input_264;
    input [44:0] input_265;
    input [44:0] input_266;
    input [44:0] input_267;
    input [44:0] input_268;
    input [44:0] input_269;
    input [44:0] input_270;
    input [44:0] input_271;
    input [44:0] input_272;
    input [44:0] input_273;
    input [44:0] input_274;
    input [44:0] input_275;
    input [44:0] input_276;
    input [44:0] input_277;
    input [44:0] input_278;
    input [44:0] input_279;
    input [44:0] input_280;
    input [44:0] input_281;
    input [44:0] input_282;
    input [44:0] input_283;
    input [44:0] input_284;
    input [44:0] input_285;
    input [44:0] input_286;
    input [44:0] input_287;
    input [44:0] input_288;
    input [44:0] input_289;
    input [44:0] input_290;
    input [44:0] input_291;
    input [44:0] input_292;
    input [44:0] input_293;
    input [44:0] input_294;
    input [44:0] input_295;
    input [44:0] input_296;
    input [44:0] input_297;
    input [44:0] input_298;
    input [44:0] input_299;
    input [44:0] input_300;
    input [44:0] input_301;
    input [44:0] input_302;
    input [44:0] input_303;
    input [44:0] input_304;
    input [44:0] input_305;
    input [44:0] input_306;
    input [44:0] input_307;
    input [44:0] input_308;
    input [44:0] input_309;
    input [44:0] input_310;
    input [44:0] input_311;
    input [44:0] input_312;
    input [44:0] input_313;
    input [44:0] input_314;
    input [44:0] input_315;
    input [44:0] input_316;
    input [44:0] input_317;
    input [44:0] input_318;
    input [44:0] input_319;
    input [44:0] input_320;
    input [44:0] input_321;
    input [44:0] input_322;
    input [44:0] input_323;
    input [8:0] sel;
    reg [44:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      default : begin
        result = input_323;
      end
    endcase
    MUX_v_45_324_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [54:0] MUX_v_55_2_2;
    input [54:0] input_0;
    input [54:0] input_1;
    input [0:0] sel;
    reg [54:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_55_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] conv_s2s_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_9_17 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_17 = {{8{vector[8]}}, vector};
  end
  endfunction


  function automatic [57:0] conv_s2s_47_58 ;
    input [46:0]  vector ;
  begin
    conv_s2s_47_58 = {{11{vector[46]}}, vector};
  end
  endfunction


  function automatic [57:0] conv_s2s_57_58 ;
    input [56:0]  vector ;
  begin
    conv_s2s_57_58 = {vector[56], vector};
  end
  endfunction


  function automatic [48:0] conv_s2u_47_49 ;
    input [46:0]  vector ;
  begin
    conv_s2u_47_49 = {{2{vector[46]}}, vector};
  end
  endfunction


  function automatic [48:0] conv_s2u_48_49 ;
    input [47:0]  vector ;
  begin
    conv_s2u_48_49 = {vector[47], vector};
  end
  endfunction


  function automatic [63:0] conv_s2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_s2u_64_64 = vector;
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [48:0] conv_u2s_1_49 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_49 = {{48{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_2_5 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_5 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_3_11 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_11 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_5_13 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_13 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_8_14 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_14 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_11_11 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_11 = vector;
  end
  endfunction


  function automatic [15:0] conv_u2u_11_16 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_16 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_13_13 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_13 = vector;
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store_core
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store_core (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_outputs_rsc_req_vz,
      plm_outputs_rsc_rls_lz, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy,
      dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, done_rsc_rdy,
      done_rsc_vld, plm_outputs_rsci_q_d, plm_outputs_rsci_radr_d, plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  input plm_outputs_rsc_req_vz;
  output plm_outputs_rsc_rls_lz;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;
  input [31:0] plm_outputs_rsci_q_d;
  output [13:0] plm_outputs_rsci_radr_d;
  output plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire core_wen;
  wire conf_info_rsci_bawt;
  wire core_wten;
  wire conf_info_rsci_wen_comp;
  wire [63:0] conf_info_rsci_idat_mxwt;
  wire plm_outputs_rsci_bawt;
  wire [31:0] plm_outputs_rsci_q_d_mxwt;
  wire dma_write_ctrl_rsci_bawt;
  wire dma_write_ctrl_rsci_wen_comp;
  wire dma_write_chnl_rsci_bawt;
  wire dma_write_chnl_rsci_wen_comp;
  wire done_rsci_bawt;
  wire done_rsci_wen_comp;
  wire plm_outputs_rsc_rls_obj_bawt;
  wire plm_outputs_rsc_req_obj_bawt;
  reg plm_outputs_rsc_req_obj_iswt0;
  wire plm_outputs_rsc_req_obj_wen_comp;
  reg [15:0] dma_write_ctrl_rsci_idat_47_32;
  reg [15:0] dma_write_ctrl_rsci_idat_15_0;
  reg [31:0] dma_write_chnl_rsci_idat_31_0;
  wire [1:0] fsm_output;
  wire [8:0] operator_8_false_1_acc_tmp;
  wire [9:0] nl_operator_8_false_1_acc_tmp;
  wire [16:0] operator_16_false_acc_tmp;
  wire [17:0] nl_operator_16_false_acc_tmp;
  wire STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_tmp;
  wire or_tmp_8;
  wire mux_tmp;
  wire mux_tmp_1;
  wire and_tmp_2;
  wire mux_tmp_33;
  wire nand_tmp_11;
  wire nand_tmp_12;
  wire mux_tmp_36;
  wire and_dcpl_5;
  wire or_dcpl_3;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire or_dcpl_4;
  wire or_dcpl_8;
  wire and_dcpl_18;
  wire and_dcpl_24;
  wire and_dcpl_26;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_36;
  wire and_dcpl_37;
  wire and_dcpl_44;
  wire and_dcpl_49;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire and_dcpl_62;
  wire and_dcpl_68;
  wire or_tmp_88;
  wire main_stage_en_5;
  wire [4:0] STORE_BATCH_LOOP_b_4_0_sva_2;
  wire [5:0] nl_STORE_BATCH_LOOP_b_4_0_sva_2;
  wire [3:0] STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1;
  wire [13:0] STORE_INNER_LOOP_i_13_0_lpi_1_dfm_mx0w0;
  reg STORE_BATCH_LOOP_asn_itm;
  reg exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1;
  reg main_stage_v_1;
  reg exit_STORE_INNER_LOOP_lpi_1_dfm_st_2;
  reg main_stage_v_2;
  reg exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4;
  reg main_stage_v_4;
  reg exitL_exit_STORE_BATCH_LOOP_sva;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2;
  reg exit_STORE_INNER_LOOP_lpi_1_dfm;
  reg exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_2;
  reg exit_STORE_INNER_LOOP_lpi_1_dfm_st_1;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_3;
  reg exit_STORE_BATCH_LOOP_sva_2;
  reg reg_conf_info_rsci_iswt0_cse;
  wire STORE_BATCH_LOOP_and_1_cse;
  reg reg_plm_outputs_rsc_rls_obj_ld_core_psct_cse;
  reg reg_done_rsci_ivld_core_psct_cse;
  reg reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  reg reg_dma_write_ctrl_rsci_ivld_core_psct_cse;
  reg reg_plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse;
  wire STORE_BATCH_LOOP_and_cse;
  wire nand_69_cse;
  wire or_171_cse;
  wire STORE_INNER_LOOP_and_cse;
  wire nor_41_cse;
  wire or_176_cse;
  wire or_183_cse;
  wire or_56_cse;
  wire and_157_cse;
  wire and_171_cse;
  wire and_163_cse;
  wire or_93_cse;
  reg [13:0] plm_outputs_rsci_radr_d_reg;
  wire [13:0] STORE_INNER_LOOP_i_mux_rmff;
  wire plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire [10:0] z_out;
  wire [10:0] z_out_1;
  wire [9:0] z_out_2;
  reg [13:0] STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1;
  reg [15:0] ac_int_cctor_8_lpi_1_dfm_1;
  reg [15:0] ac_int_cctor_8_lpi_1_dfm_2;
  reg [13:0] STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1_1;
  reg [15:0] STORE_BATCH_LOOP_acc_itm_1;
  reg [15:0] STORE_BATCH_LOOP_acc_itm_2;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2;
  reg [3:0] STORE_BATCH_LOOP_b_4_0_lpi_1_3_0;
  reg [7:0] conf_info_crt_lpi_1_dfm_231_224;
  reg [7:0] conf_info_crt_lpi_1_dfm_199_192;
  reg [7:0] conf_info_crt_lpi_1_dfm_167_160;
  reg [7:0] conf_info_crt_lpi_1_dfm_135_128;
  reg [7:0] conf_info_crt_lpi_1_dfm_103_96;
  reg [7:0] conf_info_crt_lpi_1_dfm_71_64;
  wire plm_outputs_rsc_req_obj_iswt0_mx0c1;
  wire [7:0] conf_info_crt_lpi_1_dfm_231_224_mx0;
  wire exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
  wire [13:0] STORE_INNER_LOOP_i_13_0_sva_1_mx0w0;
  wire [14:0] nl_STORE_INNER_LOOP_i_13_0_sva_1_mx0w0;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_4_mx0c1;
  wire [7:0] conf_info_crt_lpi_1_dfm_199_192_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_167_160_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_135_128_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_103_96_mx0;
  wire [7:0] conf_info_crt_lpi_1_dfm_71_64_mx0;
  wire [15:0] ac_int_cctor_8_sva_1;
  wire [23:0] nl_ac_int_cctor_8_sva_1;
  wire [7:0] pad_sva_1;
  wire signed [16:0] nl_pad_sva_1;
  wire unequal_tmp_1;
  wire [16:0] pad_acc_psp_sva_1;
  wire [17:0] nl_pad_acc_psp_sva_1;
  wire [15:0] ac_int_cctor_8_lpi_1_dfm_mx0;
  wire STORE_BATCH_LOOP_and_12_rgt;
  wire and_193_cse;
  wire STORE_INNER_LOOP_and_7_cse;
  wire STORE_BATCH_LOOP_and_13_cse;
  wire STORE_BATCH_LOOP_b_and_itm;
  wire operator_16_false_acc_itm_7_1;
  wire [1:0] if_if_and_cse;
  wire if_if_nand_2_cse;

  wire[0:0] mux_54_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] nor_47_nl;
  wire[0:0] and_101_nl;
  wire[15:0] STORE_BATCH_LOOP_acc_nl;
  wire[16:0] nl_STORE_BATCH_LOOP_acc_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_nl;
  wire[15:0] STORE_BATCH_LOOP_acc_1_nl;
  wire[16:0] nl_STORE_BATCH_LOOP_acc_1_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_1_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_1_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_2_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_3_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_3_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_4_nl;
  wire[23:0] nl_STORE_BATCH_LOOP_mul_4_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_5_nl;
  wire[15:0] STORE_BATCH_LOOP_mul_6_nl;
  wire[19:0] nl_STORE_BATCH_LOOP_mul_6_nl;
  wire[0:0] STORE_BATCH_LOOP_mux_3_nl;
  wire[0:0] STORE_INNER_LOOP_not_3_nl;
  wire[15:0] mul_1_nl;
  wire[7:0] mux_17_nl;
  wire[7:0] operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_acc_nl;
  wire[0:0] operator_42_true_and_nl;
  wire[7:0] mux_18_nl;
  wire[7:0] operator_43_true_1_acc_nl;
  wire[8:0] nl_operator_43_true_1_acc_nl;
  wire[0:0] operator_42_true_1_and_nl;
  wire[7:0] operator_43_true_operator_43_true_acc_nl;
  wire[8:0] nl_operator_43_true_operator_43_true_acc_nl;
  wire[0:0] operator_43_true_and_nl;
  wire[8:0] pad_acc_2_nl;
  wire[9:0] nl_pad_acc_2_nl;
  wire[16:0] pad_mul_nl;
  wire signed [17:0] nl_pad_mul_nl;
  wire[8:0] operator_8_false_acc_nl;
  wire[9:0] nl_operator_8_false_acc_nl;
  wire[0:0] STORE_BATCH_LOOP_not_18_nl;
  wire[7:0] operator_16_false_acc_nl;
  wire[8:0] nl_operator_16_false_acc_nl;
  wire[0:0] STORE_BATCH_LOOP_STORE_BATCH_LOOP_nor_nl;
  wire[0:0] STORE_BATCH_LOOP_and_11_nl;
  wire[0:0] and_nl;
  wire[0:0] and_10_nl;
  wire[0:0] nor_48_nl;
  wire[0:0] and_34_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] and_35_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] nor_44_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] or_142_nl;
  wire[11:0] acc_nl;
  wire[12:0] nl_acc_nl;
  wire[11:0] acc_1_nl;
  wire[12:0] nl_acc_1_nl;
  wire[10:0] acc_2_nl;
  wire[11:0] nl_acc_2_nl;
  wire[0:0] if_if_and_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_store_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg;
  assign nl_store_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg = conf_info_rsci_bawt
      & STORE_BATCH_LOOP_asn_itm & and_tmp_2 & (fsm_output[1]);
  wire [0:0] nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_oswt_unreg;
  assign nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_oswt_unreg =
      or_tmp_8 & dma_write_chnl_rsci_bawt & dma_write_ctrl_rsci_bawt & exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3
      & reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  wire [66:0] nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat;
  assign nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat = {19'b0110000000000000000
      , dma_write_ctrl_rsci_idat_47_32 , 16'b0000000000000000 , dma_write_ctrl_rsci_idat_15_0};
  wire [63:0] nl_store_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat;
  assign nl_store_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat = {32'b11011110101011011011111011101111
      , dma_write_chnl_rsci_idat_31_0};
  wire [0:0] nl_store_core_plm_outputs_rsc_rls_obj_inst_plm_outputs_rsc_rls_obj_oswt_unreg;
  assign nl_store_core_plm_outputs_rsc_rls_obj_inst_plm_outputs_rsc_rls_obj_oswt_unreg
      = mux_tmp & plm_outputs_rsci_bawt & plm_outputs_rsc_rls_obj_bawt & exit_STORE_INNER_LOOP_lpi_1_dfm_st_2
      & main_stage_v_2;
  wire [0:0] nl_store_core_plm_outputs_rsc_req_obj_inst_plm_outputs_rsc_req_obj_oswt_unreg;
  assign nl_store_core_plm_outputs_rsc_req_obj_inst_plm_outputs_rsc_req_obj_oswt_unreg
      = mux_tmp_1 & and_171_cse;
  esp_acc_conv2d_cxx_catapult_store_core_conf_info_rsci store_core_conf_info_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .core_wen(core_wen),
      .conf_info_rsci_oswt_unreg(nl_store_core_conf_info_rsci_inst_conf_info_rsci_oswt_unreg[0:0]),
      .conf_info_rsci_bawt(conf_info_rsci_bawt),
      .conf_info_rsci_iswt0(reg_conf_info_rsci_iswt0_cse),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .conf_info_rsci_idat_mxwt(conf_info_rsci_idat_mxwt)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsci_1 store_core_plm_outputs_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsci_q_d(plm_outputs_rsci_q_d),
      .plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsci_oswt_unreg(and_dcpl_33),
      .plm_outputs_rsci_bawt(plm_outputs_rsci_bawt),
      .plm_outputs_rsci_iswt0(reg_plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse),
      .plm_outputs_rsci_q_d_mxwt(plm_outputs_rsci_q_d_mxwt),
      .plm_outputs_rsci_iswt0_pff(and_dcpl_49)
    );
  esp_acc_conv2d_cxx_catapult_store_core_dma_write_ctrl_rsci store_core_dma_write_ctrl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .core_wen(core_wen),
      .dma_write_ctrl_rsci_oswt_unreg(nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_oswt_unreg[0:0]),
      .dma_write_ctrl_rsci_bawt(dma_write_ctrl_rsci_bawt),
      .dma_write_ctrl_rsci_iswt0(reg_dma_write_ctrl_rsci_ivld_core_psct_cse),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_ctrl_rsci_idat(nl_store_core_dma_write_ctrl_rsci_inst_dma_write_ctrl_rsci_idat[66:0])
    );
  esp_acc_conv2d_cxx_catapult_store_core_dma_write_chnl_rsci store_core_dma_write_chnl_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .core_wen(core_wen),
      .dma_write_chnl_rsci_oswt_unreg(and_dcpl_37),
      .dma_write_chnl_rsci_bawt(dma_write_chnl_rsci_bawt),
      .dma_write_chnl_rsci_iswt0(reg_dma_write_chnl_rsci_ivld_core_psct_cse),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .dma_write_chnl_rsci_idat(nl_store_core_dma_write_chnl_rsci_inst_dma_write_chnl_rsci_idat[63:0])
    );
  esp_acc_conv2d_cxx_catapult_store_core_done_rsci store_core_done_rsci_inst (
      .clk(clk),
      .rst(rst),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .core_wen(core_wen),
      .done_rsci_oswt_unreg(and_dcpl_29),
      .done_rsci_bawt(done_rsci_bawt),
      .done_rsci_iswt0(reg_done_rsci_ivld_core_psct_cse),
      .done_rsci_wen_comp(done_rsci_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_rls_obj store_core_plm_outputs_rsc_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_rls_lz(plm_outputs_rsc_rls_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .plm_outputs_rsc_rls_obj_oswt_unreg(nl_store_core_plm_outputs_rsc_rls_obj_inst_plm_outputs_rsc_rls_obj_oswt_unreg[0:0]),
      .plm_outputs_rsc_rls_obj_bawt(plm_outputs_rsc_rls_obj_bawt),
      .plm_outputs_rsc_rls_obj_iswt0(reg_plm_outputs_rsc_rls_obj_ld_core_psct_cse)
    );
  esp_acc_conv2d_cxx_catapult_store_core_plm_outputs_rsc_req_obj store_core_plm_outputs_rsc_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_req_vz(plm_outputs_rsc_req_vz),
      .core_wen(core_wen),
      .plm_outputs_rsc_req_obj_oswt_unreg(nl_store_core_plm_outputs_rsc_req_obj_inst_plm_outputs_rsc_req_obj_oswt_unreg[0:0]),
      .plm_outputs_rsc_req_obj_bawt(plm_outputs_rsc_req_obj_bawt),
      .plm_outputs_rsc_req_obj_iswt0(plm_outputs_rsc_req_obj_iswt0),
      .plm_outputs_rsc_req_obj_wen_comp(plm_outputs_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_store_core_staller store_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .conf_info_rsci_wen_comp(conf_info_rsci_wen_comp),
      .dma_write_ctrl_rsci_wen_comp(dma_write_ctrl_rsci_wen_comp),
      .dma_write_chnl_rsci_wen_comp(dma_write_chnl_rsci_wen_comp),
      .done_rsci_wen_comp(done_rsci_wen_comp),
      .plm_outputs_rsc_req_obj_wen_comp(plm_outputs_rsc_req_obj_wen_comp)
    );
  esp_acc_conv2d_cxx_catapult_store_core_core_fsm store_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_163_cse = or_171_cse & operator_16_false_acc_itm_7_1;
  assign or_93_cse = nor_41_cse | (STORE_BATCH_LOOP_b_4_0_sva_2[4]);
  assign STORE_BATCH_LOOP_and_cse = core_wen & (~((~ mux_tmp_33) | (fsm_output[0])));
  assign STORE_INNER_LOOP_and_cse = core_wen & (~(or_dcpl_4 | or_dcpl_3));
  assign STORE_BATCH_LOOP_and_1_cse = core_wen & (~(or_dcpl_4 | or_dcpl_8));
  assign STORE_INNER_LOOP_i_mux_rmff = MUX_v_14_2_2(STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1_1,
      plm_outputs_rsci_radr_d_reg, or_dcpl_23);
  assign or_171_cse = (operator_16_false_acc_tmp[16]) | (~((STORE_INNER_LOOP_i_13_0_lpi_1_dfm_mx0w0
      == (operator_16_false_acc_tmp[13:0])) & (operator_16_false_acc_tmp[15:14]==2'b00)));
  assign nand_69_cse = ~(or_171_cse & operator_16_false_acc_itm_7_1);
  assign STORE_BATCH_LOOP_b_and_itm = core_wen & mux_tmp_33;
  assign nor_41_cse = ~((~((STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1 == (operator_8_false_1_acc_tmp[3:0]))
      & (operator_8_false_1_acc_tmp[7:4]==4'b0000))) | (operator_8_false_1_acc_tmp[8]));
  assign STORE_BATCH_LOOP_and_12_rgt = (~ main_stage_v_1) & and_tmp_2 & (~ exitL_exit_STORE_BATCH_LOOP_sva);
  assign STORE_INNER_LOOP_and_7_cse = core_wen & and_tmp_2;
  assign STORE_BATCH_LOOP_and_13_cse = core_wen & (~ or_dcpl_22);
  assign or_176_cse = (~ exit_STORE_INNER_LOOP_lpi_1_dfm_st_2) | plm_outputs_rsc_rls_obj_bawt;
  assign and_157_cse = or_183_cse & dma_write_chnl_rsci_bawt;
  assign conf_info_crt_lpi_1_dfm_231_224_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_231_224,
      (conf_info_rsci_idat_mxwt[63:56]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign STORE_BATCH_LOOP_mux_3_nl = MUX_s_1_2_2(nor_41_cse, exit_STORE_BATCH_LOOP_sva_2,
      and_163_cse);
  assign exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0 = ((STORE_BATCH_LOOP_b_4_0_sva_2[4])
      | STORE_BATCH_LOOP_mux_3_nl) & nand_69_cse;
  assign nl_STORE_INNER_LOOP_i_13_0_sva_1_mx0w0 = STORE_INNER_LOOP_i_13_0_lpi_1_dfm_mx0w0
      + 14'b00000000000001;
  assign STORE_INNER_LOOP_i_13_0_sva_1_mx0w0 = nl_STORE_INNER_LOOP_i_13_0_sva_1_mx0w0[13:0];
  assign STORE_INNER_LOOP_not_3_nl = ~ STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_tmp;
  assign STORE_INNER_LOOP_i_13_0_lpi_1_dfm_mx0w0 = MUX_v_14_2_2(14'b00000000000000,
      STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1, STORE_INNER_LOOP_not_3_nl);
  assign STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_tmp = exit_STORE_INNER_LOOP_lpi_1_dfm
      | exit_STORE_BATCH_LOOP_lpi_1_dfm_2 | exitL_exit_STORE_BATCH_LOOP_sva;
  assign conf_info_crt_lpi_1_dfm_199_192_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_199_192,
      (conf_info_rsci_idat_mxwt[55:48]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_167_160_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_167_160,
      (conf_info_rsci_idat_mxwt[47:40]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_135_128_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_135_128,
      (conf_info_rsci_idat_mxwt[39:32]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_103_96_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_103_96,
      (conf_info_rsci_idat_mxwt[31:24]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign conf_info_crt_lpi_1_dfm_71_64_mx0 = MUX_v_8_2_2(conf_info_crt_lpi_1_dfm_71_64,
      (conf_info_rsci_idat_mxwt[23:16]), exitL_exit_STORE_BATCH_LOOP_sva);
  assign operator_42_true_and_nl = (z_out_1[10]) & (z_out_1[0]);
  assign nl_operator_43_true_acc_nl = (z_out_1[8:1]) + conv_u2s_1_8(operator_42_true_and_nl)
      + 8'b00000001;
  assign operator_43_true_acc_nl = nl_operator_43_true_acc_nl[7:0];
  assign mux_17_nl = MUX_v_8_2_2((z_out_1[7:0]), operator_43_true_acc_nl, unequal_tmp_1);
  assign operator_42_true_1_and_nl = (z_out[10]) & (z_out[0]);
  assign nl_operator_43_true_1_acc_nl = (z_out[8:1]) + conv_u2s_1_8(operator_42_true_1_and_nl)
      + 8'b00000001;
  assign operator_43_true_1_acc_nl = nl_operator_43_true_1_acc_nl[7:0];
  assign mux_18_nl = MUX_v_8_2_2((z_out[7:0]), operator_43_true_1_acc_nl, unequal_tmp_1);
  assign mul_1_nl = conv_u2u_16_16(mux_17_nl * mux_18_nl);
  assign nl_ac_int_cctor_8_sva_1 = mul_1_nl * (conf_info_rsci_idat_mxwt[23:16]);
  assign ac_int_cctor_8_sva_1 = nl_ac_int_cctor_8_sva_1[15:0];
  assign operator_43_true_and_nl = (pad_acc_psp_sva_1[16]) & (pad_acc_psp_sva_1[0]);
  assign nl_operator_43_true_operator_43_true_acc_nl = (pad_acc_psp_sva_1[8:1]) +
      conv_u2s_1_8(operator_43_true_and_nl);
  assign operator_43_true_operator_43_true_acc_nl = nl_operator_43_true_operator_43_true_acc_nl[7:0];
  assign nl_pad_sva_1 = $signed(operator_43_true_operator_43_true_acc_nl) * $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[15:8]));
  assign pad_sva_1 = nl_pad_sva_1[7:0];
  assign unequal_tmp_1 = ~((conf_info_rsci_idat_mxwt[7:0]==8'b00000001));
  assign nl_pad_acc_2_nl = ({1'b1 , (~ (conf_info_rsci_idat_mxwt[55:48]))}) + conv_u2s_8_9(conf_info_rsci_idat_mxwt[31:24])
      + 9'b000000001;
  assign pad_acc_2_nl = nl_pad_acc_2_nl[8:0];
  assign nl_operator_8_false_acc_nl = conv_u2s_8_9(conf_info_rsci_idat_mxwt[55:48])
      + 9'b111111111;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[8:0];
  assign nl_pad_mul_nl = $signed(conv_u2s_8_9(conf_info_rsci_idat_mxwt[7:0])) * $signed(operator_8_false_acc_nl);
  assign pad_mul_nl = nl_pad_mul_nl[16:0];
  assign nl_pad_acc_psp_sva_1 = conv_s2s_9_17(pad_acc_2_nl) + pad_mul_nl;
  assign pad_acc_psp_sva_1 = nl_pad_acc_psp_sva_1[16:0];
  assign nl_STORE_BATCH_LOOP_b_4_0_sva_2 = conv_u2u_4_5(STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1)
      + 5'b00001;
  assign STORE_BATCH_LOOP_b_4_0_sva_2 = nl_STORE_BATCH_LOOP_b_4_0_sva_2[4:0];
  assign STORE_BATCH_LOOP_not_18_nl = ~ exitL_exit_STORE_BATCH_LOOP_sva;
  assign STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1 = MUX_v_4_2_2(4'b0000, STORE_BATCH_LOOP_b_4_0_lpi_1_3_0,
      STORE_BATCH_LOOP_not_18_nl);
  assign nl_operator_8_false_1_acc_tmp = conv_u2s_8_9(conf_info_crt_lpi_1_dfm_231_224_mx0)
      + 9'b111111111;
  assign operator_8_false_1_acc_tmp = nl_operator_8_false_1_acc_tmp[8:0];
  assign nl_operator_16_false_acc_nl = conv_u2s_7_8(STORE_INNER_LOOP_i_13_0_sva_1_mx0w0[13:7])
      + 8'b10101111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[7:0];
  assign operator_16_false_acc_itm_7_1 = readslicef_8_1_7(operator_16_false_acc_nl);
  assign nl_operator_16_false_acc_tmp = conv_u2s_16_17(ac_int_cctor_8_lpi_1_dfm_mx0)
      + 17'b11111111111111111;
  assign operator_16_false_acc_tmp = nl_operator_16_false_acc_tmp[16:0];
  assign STORE_BATCH_LOOP_STORE_BATCH_LOOP_nor_nl = ~(main_stage_v_1 | exitL_exit_STORE_BATCH_LOOP_sva);
  assign STORE_BATCH_LOOP_and_11_nl = main_stage_v_1 & (~ exitL_exit_STORE_BATCH_LOOP_sva);
  assign ac_int_cctor_8_lpi_1_dfm_mx0 = MUX1HOT_v_16_3_2(STORE_BATCH_LOOP_acc_itm_1,
      ac_int_cctor_8_lpi_1_dfm_1, ac_int_cctor_8_sva_1, {STORE_BATCH_LOOP_STORE_BATCH_LOOP_nor_nl
      , STORE_BATCH_LOOP_and_11_nl , exitL_exit_STORE_BATCH_LOOP_sva});
  assign main_stage_en_5 = ((~ STORE_BATCH_LOOP_asn_itm) | conf_info_rsci_bawt) &
      (plm_outputs_rsc_req_obj_bawt | (~(exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1
      & main_stage_v_1))) & (plm_outputs_rsci_bawt | (~ main_stage_v_2)) & (plm_outputs_rsc_rls_obj_bawt
      | (~(exit_STORE_INNER_LOOP_lpi_1_dfm_st_2 & main_stage_v_2))) & (dma_write_ctrl_rsci_bawt
      | (~(exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3 & reg_dma_write_chnl_rsci_ivld_core_psct_cse)))
      & (dma_write_chnl_rsci_bawt | (~ reg_dma_write_chnl_rsci_ivld_core_psct_cse))
      & (done_rsci_bawt | (~(exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4 & main_stage_v_4)));
  assign or_tmp_8 = (~ main_stage_v_4) | done_rsci_bawt | (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4);
  assign or_183_cse = (~ exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3) | dma_write_ctrl_rsci_bawt;
  assign and_nl = or_183_cse & dma_write_chnl_rsci_bawt & or_tmp_8;
  assign mux_tmp = MUX_s_1_2_2(or_tmp_8, and_nl, reg_dma_write_chnl_rsci_ivld_core_psct_cse);
  assign and_10_nl = or_176_cse & plm_outputs_rsci_bawt & mux_tmp;
  assign mux_tmp_1 = MUX_s_1_2_2(mux_tmp, and_10_nl, main_stage_v_2);
  assign and_tmp_2 = ((~ main_stage_v_1) | (~ exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1)
      | plm_outputs_rsc_req_obj_bawt) & mux_tmp_1;
  assign or_56_cse = (~ exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1) | plm_outputs_rsc_req_obj_bawt;
  assign and_171_cse = main_stage_v_1 & exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1
      & plm_outputs_rsc_req_obj_bawt;
  assign nor_48_nl = ~(STORE_BATCH_LOOP_asn_itm | (~ and_tmp_2));
  assign mux_tmp_33 = MUX_s_1_2_2(nor_48_nl, and_tmp_2, conf_info_rsci_bawt);
  assign nand_tmp_11 = ~(exitL_exit_STORE_BATCH_LOOP_sva & (~ mux_tmp_33));
  assign nand_tmp_12 = ~(reg_dma_write_chnl_rsci_ivld_core_psct_cse & (~ and_157_cse));
  assign and_34_nl = or_176_cse & plm_outputs_rsci_bawt & nand_tmp_12;
  assign mux_tmp_36 = MUX_s_1_2_2(nand_tmp_12, and_34_nl, main_stage_v_2);
  assign and_dcpl_5 = (~ plm_outputs_rsc_rls_obj_bawt) & exit_STORE_INNER_LOOP_lpi_1_dfm_st_2;
  assign or_dcpl_3 = and_dcpl_5 | (~ plm_outputs_rsci_bawt) | (~ main_stage_v_2);
  assign and_dcpl_7 = (~ done_rsci_bawt) & exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4
      & main_stage_v_4;
  assign and_dcpl_8 = (~ and_157_cse) & reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  assign or_dcpl_4 = and_dcpl_8 | and_dcpl_7;
  assign or_dcpl_8 = and_dcpl_5 | (~ plm_outputs_rsci_bawt) | (~(main_stage_v_2 &
      exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_2));
  assign and_dcpl_18 = mux_tmp_1 & or_56_cse;
  assign and_dcpl_24 = dma_write_chnl_rsci_bawt & reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  assign and_dcpl_26 = or_tmp_8 & or_183_cse;
  assign and_dcpl_29 = done_rsci_bawt & exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4 &
      main_stage_v_4;
  assign and_dcpl_30 = (~(and_157_cse & reg_dma_write_chnl_rsci_ivld_core_psct_cse
      & exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_3)) & and_dcpl_29;
  assign and_dcpl_31 = plm_outputs_rsci_bawt & main_stage_v_2;
  assign and_dcpl_32 = mux_tmp & or_176_cse;
  assign and_dcpl_33 = and_dcpl_32 & and_dcpl_31;
  assign and_dcpl_36 = or_dcpl_3 & or_tmp_8 & or_183_cse & and_dcpl_24;
  assign and_dcpl_37 = and_dcpl_26 & and_dcpl_24;
  assign and_dcpl_44 = or_dcpl_8 & or_tmp_8 & dma_write_chnl_rsci_bawt & dma_write_ctrl_rsci_bawt
      & exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3 & reg_dma_write_chnl_rsci_ivld_core_psct_cse;
  assign and_dcpl_49 = and_dcpl_18 & main_stage_v_1;
  assign or_dcpl_22 = (~ mux_tmp_36) | and_dcpl_7;
  assign or_dcpl_23 = or_dcpl_22 | (~((~((~ plm_outputs_rsc_req_obj_bawt) & exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1))
      & main_stage_v_1));
  assign and_dcpl_62 = and_dcpl_18 & main_stage_v_1 & STORE_BATCH_LOOP_asn_itm &
      (~ conf_info_rsci_bawt);
  assign and_dcpl_68 = (~ dma_write_ctrl_rsci_bawt) & exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3;
  assign and_35_nl = or_171_cse & operator_16_false_acc_itm_7_1 & mux_tmp_36;
  assign mux_56_nl = MUX_s_1_2_2(mux_tmp_36, and_35_nl, or_93_cse);
  assign mux_57_nl = MUX_s_1_2_2(mux_tmp_36, mux_56_nl, main_stage_en_5);
  assign or_tmp_88 = mux_57_nl & or_tmp_8 & (or_56_cse | (~ main_stage_v_1)) & STORE_BATCH_LOOP_asn_itm
      & conf_info_rsci_bawt & (fsm_output[1]);
  assign nor_44_nl = ~(conf_info_rsci_bawt | (~(STORE_BATCH_LOOP_asn_itm & mux_tmp_36)));
  assign mux_62_nl = MUX_s_1_2_2(mux_tmp_36, nor_44_nl, STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_tmp);
  assign plm_outputs_rsc_req_obj_iswt0_mx0c1 = mux_62_nl & or_tmp_8 & and_171_cse;
  assign or_142_nl = or_56_cse | and_dcpl_8;
  assign mux_74_nl = MUX_s_1_2_2(and_dcpl_8, or_142_nl, main_stage_v_1);
  assign main_stage_v_2_mx0c1 = (~ mux_74_nl) & or_tmp_8 & or_176_cse & and_dcpl_31;
  assign main_stage_v_4_mx0c1 = (and_dcpl_68 | (~ dma_write_chnl_rsci_bawt) | (~
      reg_dma_write_chnl_rsci_ivld_core_psct_cse)) & (done_rsci_bawt | (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4))
      & main_stage_v_4;
  assign plm_outputs_rsci_radr_d = STORE_INNER_LOOP_i_mux_rmff;
  assign plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d = plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign and_193_cse = ((conf_info_rsci_idat_mxwt[7:0]!=8'b00000001)) & (fsm_output[1]);
  assign if_if_and_cse = MUX_v_2_2_2(2'b00, (z_out_2[9:8]), and_193_cse);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_conf_info_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (((~ mux_54_nl) & main_stage_en_5) | (fsm_output[0]) | or_tmp_88)
        ) begin
      reg_conf_info_rsci_iswt0_cse <= ~ or_tmp_88;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exitL_exit_STORE_BATCH_LOOP_sva <= 1'b1;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2 <= 1'b0;
      exit_STORE_INNER_LOOP_lpi_1_dfm <= 1'b0;
      exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1 <= 1'b0;
    end
    else if ( STORE_BATCH_LOOP_and_cse ) begin
      exitL_exit_STORE_BATCH_LOOP_sva <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
      exit_STORE_INNER_LOOP_lpi_1_dfm <= nand_69_cse;
      exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1 <= STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_tmp;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_rsci_idat_31_0 <= 32'b00000000000000000000000000000000;
      exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3 <= 1'b0;
    end
    else if ( STORE_INNER_LOOP_and_cse ) begin
      dma_write_chnl_rsci_idat_31_0 <= plm_outputs_rsci_q_d_mxwt;
      exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_3 <= exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_rsci_idat_15_0 <= 16'b0000000000000000;
      dma_write_ctrl_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( STORE_BATCH_LOOP_and_1_cse ) begin
      dma_write_ctrl_rsci_idat_15_0 <= STORE_BATCH_LOOP_acc_itm_2;
      dma_write_ctrl_rsci_idat_47_32 <= ac_int_cctor_8_lpi_1_dfm_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_outputs_rsc_req_obj_iswt0 <= 1'b0;
    end
    else if ( core_wen & ((mux_tmp_33 & STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_tmp
        & (fsm_output[1])) | (mux_tmp_33 & (exit_STORE_BATCH_LOOP_lpi_1_dfm_2 | exit_STORE_INNER_LOOP_lpi_1_dfm)
        & (~ exitL_exit_STORE_BATCH_LOOP_sva)) | plm_outputs_rsc_req_obj_iswt0_mx0c1)
        ) begin
      plm_outputs_rsc_req_obj_iswt0 <= ~ plm_outputs_rsc_req_obj_iswt0_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_plm_outputs_rsc_rls_obj_ld_core_psct_cse <= 1'b0;
      reg_plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= 1'b0;
      plm_outputs_rsci_radr_d_reg <= 14'b00000000000000;
      conf_info_crt_lpi_1_dfm_231_224 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_199_192 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_167_160 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_135_128 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_103_96 <= 8'b00000000;
      conf_info_crt_lpi_1_dfm_71_64 <= 8'b00000000;
    end
    else if ( core_wen ) begin
      reg_plm_outputs_rsc_rls_obj_ld_core_psct_cse <= and_dcpl_18 & main_stage_v_1
          & exit_STORE_INNER_LOOP_lpi_1_dfm_st_1;
      reg_plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d_core_psct_cse <= and_dcpl_49;
      plm_outputs_rsci_radr_d_reg <= STORE_INNER_LOOP_i_mux_rmff;
      conf_info_crt_lpi_1_dfm_231_224 <= conf_info_crt_lpi_1_dfm_231_224_mx0;
      conf_info_crt_lpi_1_dfm_199_192 <= conf_info_crt_lpi_1_dfm_199_192_mx0;
      conf_info_crt_lpi_1_dfm_167_160 <= conf_info_crt_lpi_1_dfm_167_160_mx0;
      conf_info_crt_lpi_1_dfm_135_128 <= conf_info_crt_lpi_1_dfm_135_128_mx0;
      conf_info_crt_lpi_1_dfm_103_96 <= conf_info_crt_lpi_1_dfm_103_96_mx0;
      conf_info_crt_lpi_1_dfm_71_64 <= conf_info_crt_lpi_1_dfm_71_64_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_done_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_26 & and_dcpl_24 & exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_3)
        | and_dcpl_30) ) begin
      reg_done_rsci_ivld_core_psct_cse <= ~ and_dcpl_30;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_write_chnl_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_33 | and_dcpl_36) ) begin
      reg_dma_write_chnl_rsci_ivld_core_psct_cse <= ~ and_dcpl_36;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_write_ctrl_rsci_ivld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_32 & and_dcpl_31 & exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_2)
        | and_dcpl_44) ) begin
      reg_dma_write_ctrl_rsci_ivld_core_psct_cse <= ~ and_dcpl_44;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_asn_itm <= 1'b1;
    end
    else if ( core_wen & ((main_stage_en_5 & (fsm_output[1])) | ((~ STORE_BATCH_LOOP_asn_itm)
        & main_stage_en_5)) ) begin
      STORE_BATCH_LOOP_asn_itm <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~((~ mux_tmp_33) | and_163_cse | (fsm_output[0]))) ) begin
      exit_STORE_BATCH_LOOP_sva_2 <= nor_41_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_b_4_0_lpi_1_3_0 <= 4'b0000;
      STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1 <= 14'b00000000000000;
    end
    else if ( STORE_BATCH_LOOP_b_and_itm ) begin
      STORE_BATCH_LOOP_b_4_0_lpi_1_3_0 <= MUX_v_4_2_2((STORE_BATCH_LOOP_b_4_0_sva_2[3:0]),
          STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1, and_101_nl);
      STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1 <= STORE_INNER_LOOP_i_13_0_sva_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & ((mux_tmp_33 & (fsm_output[1])) | and_dcpl_62) ) begin
      main_stage_v_1 <= ~ and_dcpl_62;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      ac_int_cctor_8_lpi_1_dfm_1 <= 16'b0000000000000000;
    end
    else if ( core_wen & ((and_tmp_2 & exitL_exit_STORE_BATCH_LOOP_sva) | STORE_BATCH_LOOP_and_12_rgt)
        ) begin
      ac_int_cctor_8_lpi_1_dfm_1 <= MUX_v_16_2_2(ac_int_cctor_8_sva_1, STORE_BATCH_LOOP_acc_itm_1,
          STORE_BATCH_LOOP_and_12_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_INNER_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1_1 <= 14'b00000000000000;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1 <= 1'b0;
    end
    else if ( STORE_INNER_LOOP_and_7_cse ) begin
      exit_STORE_INNER_LOOP_lpi_1_dfm_st_1 <= nand_69_cse;
      STORE_INNER_LOOP_i_13_0_lpi_1_dfm_1_1 <= STORE_INNER_LOOP_i_13_0_lpi_1_dfm_mx0w0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_49 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_acc_itm_2 <= 16'b0000000000000000;
      ac_int_cctor_8_lpi_1_dfm_2 <= 16'b0000000000000000;
      exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2 <= 1'b0;
    end
    else if ( STORE_BATCH_LOOP_and_13_cse ) begin
      STORE_BATCH_LOOP_acc_itm_2 <= STORE_BATCH_LOOP_acc_itm_1;
      ac_int_cctor_8_lpi_1_dfm_2 <= ac_int_cctor_8_lpi_1_dfm_1;
      exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_2 <= exitL_exit_STORE_INNER_LOOP_lpi_1_dfm_st_1;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_INNER_LOOP_lpi_1_dfm_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_23) ) begin
      exit_STORE_INNER_LOOP_lpi_1_dfm_st_2 <= exit_STORE_INNER_LOOP_lpi_1_dfm_st_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_3 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_4) ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_3 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_37 | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4 <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_7 | (~ dma_write_chnl_rsci_bawt) | and_dcpl_68
        | (~ reg_dma_write_chnl_rsci_ivld_core_psct_cse))) ) begin
      exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_4 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_2_st_3;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_acc_itm_1 <= 16'b0000000000000000;
    end
    else if ( core_wen & (mux_tmp_33 | and_dcpl_62) ) begin
      STORE_BATCH_LOOP_acc_itm_1 <= MUX_v_16_2_2(STORE_BATCH_LOOP_acc_nl, ac_int_cctor_8_lpi_1_dfm_1,
          and_dcpl_62);
    end
  end
  assign nor_47_nl = ~(exitL_exit_STORE_BATCH_LOOP_sva | mux_tmp_33);
  assign mux_53_nl = MUX_s_1_2_2(nor_47_nl, nand_tmp_11, and_163_cse);
  assign mux_54_nl = MUX_s_1_2_2(nand_tmp_11, mux_53_nl, or_93_cse);
  assign and_101_nl = mux_tmp_33 & and_163_cse;
  assign STORE_BATCH_LOOP_mul_2_nl = conv_u2u_16_16(conf_info_crt_lpi_1_dfm_199_192_mx0
      * conf_info_crt_lpi_1_dfm_167_160_mx0);
  assign nl_STORE_BATCH_LOOP_mul_1_nl = STORE_BATCH_LOOP_mul_2_nl * conf_info_crt_lpi_1_dfm_135_128_mx0;
  assign STORE_BATCH_LOOP_mul_1_nl = nl_STORE_BATCH_LOOP_mul_1_nl[15:0];
  assign STORE_BATCH_LOOP_mul_5_nl = conv_u2u_16_16(conf_info_crt_lpi_1_dfm_103_96_mx0
      * conf_info_crt_lpi_1_dfm_103_96_mx0);
  assign nl_STORE_BATCH_LOOP_mul_4_nl = STORE_BATCH_LOOP_mul_5_nl * conf_info_crt_lpi_1_dfm_135_128_mx0;
  assign STORE_BATCH_LOOP_mul_4_nl = nl_STORE_BATCH_LOOP_mul_4_nl[15:0];
  assign nl_STORE_BATCH_LOOP_mul_3_nl = STORE_BATCH_LOOP_mul_4_nl * conf_info_crt_lpi_1_dfm_71_64_mx0;
  assign STORE_BATCH_LOOP_mul_3_nl = nl_STORE_BATCH_LOOP_mul_3_nl[15:0];
  assign nl_STORE_BATCH_LOOP_acc_1_nl = STORE_BATCH_LOOP_mul_1_nl + STORE_BATCH_LOOP_mul_3_nl;
  assign STORE_BATCH_LOOP_acc_1_nl = nl_STORE_BATCH_LOOP_acc_1_nl[15:0];
  assign nl_STORE_BATCH_LOOP_mul_nl = conf_info_crt_lpi_1_dfm_231_224_mx0 * STORE_BATCH_LOOP_acc_1_nl;
  assign STORE_BATCH_LOOP_mul_nl = nl_STORE_BATCH_LOOP_mul_nl[15:0];
  assign nl_STORE_BATCH_LOOP_mul_6_nl = ac_int_cctor_8_lpi_1_dfm_mx0 * STORE_BATCH_LOOP_b_4_0_lpi_1_dfm_3_0_1;
  assign STORE_BATCH_LOOP_mul_6_nl = nl_STORE_BATCH_LOOP_mul_6_nl[15:0];
  assign nl_STORE_BATCH_LOOP_acc_nl = STORE_BATCH_LOOP_mul_nl + STORE_BATCH_LOOP_mul_6_nl;
  assign STORE_BATCH_LOOP_acc_nl = nl_STORE_BATCH_LOOP_acc_nl[15:0];
  assign if_if_nand_2_cse = ~(and_193_cse & (~((conf_info_rsci_idat_mxwt[7:0]==8'b00000001)
      & (fsm_output[1]))));
  assign nl_acc_nl = conv_u2u_11_12({if_if_and_cse , (z_out_2[7:0]) , if_if_nand_2_cse})
      + conv_s2u_10_12({and_193_cse , (conf_info_rsci_idat_mxwt[47:40]) , 1'b1});
  assign acc_nl = nl_acc_nl[11:0];
  assign z_out = readslicef_12_11_1(acc_nl);
  assign nl_acc_1_nl = conv_u2u_11_12({if_if_and_cse , (z_out_2[7:0]) , if_if_nand_2_cse})
      + conv_s2u_10_12({and_193_cse , (conf_info_rsci_idat_mxwt[55:48]) , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[11:0];
  assign z_out_1 = readslicef_12_11_1(acc_1_nl);
  assign if_if_and_3_nl = (pad_sva_1[7]) & and_193_cse;
  assign nl_acc_2_nl = conv_u2u_10_11({if_if_and_3_nl , (pad_sva_1[6:0]) , 2'b01})
      + conv_u2u_9_11({(~ (conf_info_rsci_idat_mxwt[31:24])) , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[10:0];
  assign z_out_2 = readslicef_11_10_1(acc_2_nl);

  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [16:0] conv_s2s_9_17 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_17 = {{8{vector[8]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_10_12 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_12 = {{2{vector[9]}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_8 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [16:0] conv_u2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_17 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_16 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core (
  clk, rst, acc_done_rsc_vld, config_done_cns_rdy, config_done_cns_vld, load_done_cns_rdy,
      load_done_cns_vld, compute_done_cns_rdy, compute_done_cns_vld, store_done_cns_rdy,
      store_done_cns_vld
);
  input clk;
  input rst;
  output acc_done_rsc_vld;
  output config_done_cns_rdy;
  input config_done_cns_vld;
  output load_done_cns_rdy;
  input load_done_cns_vld;
  output compute_done_cns_rdy;
  input compute_done_cns_vld;
  output store_done_cns_rdy;
  input store_done_cns_vld;



  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core_core conv2d_cxx_catapult_core_core_inst
      (
      .clk(clk),
      .rst(rst),
      .acc_done_rsc_vld(acc_done_rsc_vld),
      .config_done_cns_rdy(config_done_cns_rdy),
      .config_done_cns_vld(config_done_cns_vld),
      .load_done_cns_rdy(load_done_cns_rdy),
      .load_done_cns_vld(load_done_cns_vld),
      .compute_done_cns_rdy(compute_done_cns_rdy),
      .compute_done_cns_vld(compute_done_cns_vld),
      .store_done_cns_rdy(store_done_cns_rdy),
      .store_done_cns_vld(store_done_cns_vld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_config
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_config (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_conf_load_rsc_dat,
      plm_conf_load_rsc_vld, plm_conf_load_rsc_rdy, plm_conf_compute_rsc_dat, plm_conf_compute_rsc_vld,
      plm_conf_compute_rsc_rdy, plm_conf_store_rsc_dat, plm_conf_store_rsc_vld, plm_conf_store_rsc_rdy,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [255:0] plm_conf_load_rsc_dat;
  output plm_conf_load_rsc_vld;
  input plm_conf_load_rsc_rdy;
  output [255:0] plm_conf_compute_rsc_dat;
  output plm_conf_compute_rsc_vld;
  input plm_conf_compute_rsc_rdy;
  output [255:0] plm_conf_store_rsc_dat;
  output plm_conf_store_rsc_vld;
  input plm_conf_store_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;



  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_config_core config_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .plm_conf_load_rsc_dat(plm_conf_load_rsc_dat),
      .plm_conf_load_rsc_vld(plm_conf_load_rsc_vld),
      .plm_conf_load_rsc_rdy(plm_conf_load_rsc_rdy),
      .plm_conf_compute_rsc_dat(plm_conf_compute_rsc_dat),
      .plm_conf_compute_rsc_vld(plm_conf_compute_rsc_vld),
      .plm_conf_compute_rsc_rdy(plm_conf_compute_rsc_rdy),
      .plm_conf_store_rsc_dat(plm_conf_store_rsc_dat),
      .plm_conf_store_rsc_vld(plm_conf_store_rsc_vld),
      .plm_conf_store_rsc_rdy(plm_conf_store_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_load
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_load (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_inputs_rsc_wadr,
      plm_inputs_rsc_d, plm_inputs_rsc_we, plm_inputs_rsc_req_vz, plm_inputs_rsc_rls_lz,
      plm_filters_rsc_wadr, plm_filters_rsc_d, plm_filters_rsc_we, plm_filters_rsc_req_vz,
      plm_filters_rsc_rls_lz, dma_read_ctrl_rsc_dat, dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy,
      dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy, done_rsc_rdy,
      done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [13:0] plm_inputs_rsc_wadr;
  output [31:0] plm_inputs_rsc_d;
  output plm_inputs_rsc_we;
  input plm_inputs_rsc_req_vz;
  output plm_inputs_rsc_rls_lz;
  output [15:0] plm_filters_rsc_wadr;
  output [31:0] plm_filters_rsc_d;
  output plm_filters_rsc_we;
  input plm_filters_rsc_req_vz;
  output plm_filters_rsc_rls_lz;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire [31:0] plm_inputs_rsci_d_d;
  wire [13:0] plm_inputs_rsci_wadr_d;
  wire [31:0] plm_filters_rsci_d_d;
  wire [15:0] plm_filters_rsci_wadr_d;
  wire plm_inputs_rsci_we_d_iff;
  wire plm_filters_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_7_14_32_10368_10368_32_1_gen
      plm_inputs_rsci (
      .we(plm_inputs_rsc_we),
      .d(plm_inputs_rsc_d),
      .wadr(plm_inputs_rsc_wadr),
      .d_d(plm_inputs_rsci_d_d),
      .wadr_d(plm_inputs_rsci_wadr_d),
      .we_d(plm_inputs_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_inputs_rsci_we_d_iff)
    );
  esp_acc_conv2d_cxx_catapult_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_8_16_32_50176_50176_32_1_gen
      plm_filters_rsci (
      .we(plm_filters_rsc_we),
      .d(plm_filters_rsc_d),
      .wadr(plm_filters_rsc_wadr),
      .d_d(plm_filters_rsci_d_d),
      .wadr_d(plm_filters_rsci_wadr_d),
      .we_d(plm_filters_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_filters_rsci_we_d_iff)
    );
  esp_acc_conv2d_cxx_catapult_load_core load_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .plm_inputs_rsc_req_vz(plm_inputs_rsc_req_vz),
      .plm_inputs_rsc_rls_lz(plm_inputs_rsc_rls_lz),
      .plm_filters_rsc_req_vz(plm_filters_rsc_req_vz),
      .plm_filters_rsc_rls_lz(plm_filters_rsc_rls_lz),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .plm_inputs_rsci_d_d(plm_inputs_rsci_d_d),
      .plm_inputs_rsci_wadr_d(plm_inputs_rsci_wadr_d),
      .plm_filters_rsci_d_d(plm_filters_rsci_d_d),
      .plm_filters_rsci_wadr_d(plm_filters_rsci_wadr_d),
      .plm_inputs_rsci_we_d_pff(plm_inputs_rsci_we_d_iff),
      .plm_filters_rsci_we_d_pff(plm_filters_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_compute
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_compute (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_inputs_rsc_radr,
      plm_inputs_rsc_q, plm_inputs_rsc_req_vz, plm_inputs_rsc_rls_lz, plm_filters_rsc_radr,
      plm_filters_rsc_q, plm_filters_rsc_req_vz, plm_filters_rsc_rls_lz, plm_outputs_rsc_wadr,
      plm_outputs_rsc_d, plm_outputs_rsc_we, plm_outputs_rsc_req_vz, plm_outputs_rsc_rls_lz,
      done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [13:0] plm_inputs_rsc_radr;
  input [31:0] plm_inputs_rsc_q;
  input plm_inputs_rsc_req_vz;
  output plm_inputs_rsc_rls_lz;
  output [15:0] plm_filters_rsc_radr;
  input [31:0] plm_filters_rsc_q;
  input plm_filters_rsc_req_vz;
  output plm_filters_rsc_rls_lz;
  output [13:0] plm_outputs_rsc_wadr;
  output [31:0] plm_outputs_rsc_d;
  output plm_outputs_rsc_we;
  input plm_outputs_rsc_req_vz;
  output plm_outputs_rsc_rls_lz;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire [31:0] plm_inputs_rsci_q_d;
  wire [13:0] plm_inputs_rsci_radr_d;
  wire plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_filters_rsci_q_d;
  wire [15:0] plm_filters_rsci_radr_d;
  wire plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_outputs_rsci_d_d;
  wire [13:0] plm_outputs_rsci_wadr_d;
  wire plm_outputs_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_15_14_32_10368_10368_32_1_gen
      plm_inputs_rsci (
      .q(plm_inputs_rsc_q),
      .radr(plm_inputs_rsc_radr),
      .q_d(plm_inputs_rsci_q_d),
      .radr_d(plm_inputs_rsci_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_16_16_32_50176_50176_32_1_gen
      plm_filters_rsci (
      .q(plm_filters_rsc_q),
      .radr(plm_filters_rsc_radr),
      .q_d(plm_filters_rsci_q_d),
      .radr_d(plm_filters_rsci_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_conv2d_cxx_catapult_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_17_14_32_10368_10368_32_1_gen
      plm_outputs_rsci (
      .we(plm_outputs_rsc_we),
      .d(plm_outputs_rsc_d),
      .wadr(plm_outputs_rsc_wadr),
      .d_d(plm_outputs_rsci_d_d),
      .wadr_d(plm_outputs_rsci_wadr_d),
      .we_d(plm_outputs_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_outputs_rsci_we_d_iff)
    );
  esp_acc_conv2d_cxx_catapult_compute_core compute_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .plm_inputs_rsc_req_vz(plm_inputs_rsc_req_vz),
      .plm_inputs_rsc_rls_lz(plm_inputs_rsc_rls_lz),
      .plm_filters_rsc_req_vz(plm_filters_rsc_req_vz),
      .plm_filters_rsc_rls_lz(plm_filters_rsc_rls_lz),
      .plm_outputs_rsc_req_vz(plm_outputs_rsc_req_vz),
      .plm_outputs_rsc_rls_lz(plm_outputs_rsc_rls_lz),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .plm_inputs_rsci_q_d(plm_inputs_rsci_q_d),
      .plm_inputs_rsci_radr_d(plm_inputs_rsci_radr_d),
      .plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_inputs_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_filters_rsci_q_d(plm_filters_rsci_q_d),
      .plm_filters_rsci_radr_d(plm_filters_rsci_radr_d),
      .plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_filters_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_outputs_rsci_d_d(plm_outputs_rsci_d_d),
      .plm_outputs_rsci_wadr_d(plm_outputs_rsci_wadr_d),
      .plm_outputs_rsci_we_d_pff(plm_outputs_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_store
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_store (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, plm_outputs_rsc_radr,
      plm_outputs_rsc_q, plm_outputs_rsc_req_vz, plm_outputs_rsc_rls_lz, dma_write_ctrl_rsc_dat,
      dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy, dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld,
      dma_write_chnl_rsc_rdy, done_rsc_rdy, done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [13:0] plm_outputs_rsc_radr;
  input [31:0] plm_outputs_rsc_q;
  input plm_outputs_rsc_req_vz;
  output plm_outputs_rsc_rls_lz;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  input done_rsc_rdy;
  output done_rsc_vld;


  // Interconnect Declarations
  wire [31:0] plm_outputs_rsci_q_d;
  wire [13:0] plm_outputs_rsci_radr_d;
  wire plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_conv2d_cxx_catapult_store_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_24_14_32_10368_10368_32_1_gen
      plm_outputs_rsci (
      .q(plm_outputs_rsc_q),
      .radr(plm_outputs_rsc_radr),
      .q_d(plm_outputs_rsci_q_d),
      .radr_d(plm_outputs_rsci_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_conv2d_cxx_catapult_store_core store_core_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .plm_outputs_rsc_req_vz(plm_outputs_rsc_req_vz),
      .plm_outputs_rsc_rls_lz(plm_outputs_rsc_rls_lz),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy),
      .done_rsc_vld(done_rsc_vld),
      .plm_outputs_rsci_q_d(plm_outputs_rsci_q_d),
      .plm_outputs_rsci_radr_d(plm_outputs_rsci_radr_d),
      .plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d(plm_outputs_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_struct
// ------------------------------------------------------------------


module esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_struct (
  clk, rst, conf_info_rsc_dat_batch, conf_info_rsc_dat_n_w, conf_info_rsc_dat_n_h,
      conf_info_rsc_dat_n_c, conf_info_rsc_dat_kern, conf_info_rsc_dat_filt, conf_info_rsc_dat_same,
      conf_info_rsc_dat_stride, conf_info_rsc_vld, conf_info_rsc_rdy, dma_read_ctrl_rsc_dat_size,
      dma_read_ctrl_rsc_dat_length, dma_read_ctrl_rsc_dat_index, dma_read_ctrl_rsc_vld,
      dma_read_ctrl_rsc_rdy, dma_write_ctrl_rsc_dat_size, dma_write_ctrl_rsc_dat_length,
      dma_write_ctrl_rsc_dat_index, dma_write_ctrl_rsc_vld, dma_write_ctrl_rsc_rdy,
      dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy, dma_write_chnl_rsc_dat,
      dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, acc_done_rsc_vld
);
  input clk;
  input rst;
  input [31:0] conf_info_rsc_dat_batch;
  input [31:0] conf_info_rsc_dat_n_w;
  input [31:0] conf_info_rsc_dat_n_h;
  input [31:0] conf_info_rsc_dat_n_c;
  input [31:0] conf_info_rsc_dat_kern;
  input [31:0] conf_info_rsc_dat_filt;
  input [31:0] conf_info_rsc_dat_same;
  input [31:0] conf_info_rsc_dat_stride;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [2:0] dma_read_ctrl_rsc_dat_size;
  output [31:0] dma_read_ctrl_rsc_dat_length;
  output [31:0] dma_read_ctrl_rsc_dat_index;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  output [2:0] dma_write_ctrl_rsc_dat_size;
  output [31:0] dma_write_ctrl_rsc_dat_length;
  output [31:0] dma_write_ctrl_rsc_dat_index;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  output acc_done_rsc_vld;


  // Interconnect Declarations
  wire [255:0] plm_conf_load_rsc_dat_nconfig_inst;
  wire plm_conf_load_rsc_rdy_nconfig_inst;
  wire [255:0] plm_conf_compute_rsc_dat_nconfig_inst;
  wire plm_conf_compute_rsc_rdy_nconfig_inst;
  wire [255:0] plm_conf_store_rsc_dat_nconfig_inst;
  wire plm_conf_store_rsc_rdy_nconfig_inst;
  wire done_rsc_rdy_nconfig_inst;
  wire [255:0] conf_info_rsc_dat_nload_inst;
  wire conf_info_rsc_vld_nload_inst;
  wire conf_info_rsc_rdy_nload_inst;
  wire [13:0] plm_inputs_rsc_wadr_nload_inst;
  wire [31:0] plm_inputs_rsc_d_nload_inst;
  wire plm_inputs_rsc_we_nload_inst;
  wire plm_inputs_rsc_req_vz_nload_inst;
  wire [15:0] plm_filters_rsc_wadr_nload_inst;
  wire [31:0] plm_filters_rsc_d_nload_inst;
  wire plm_filters_rsc_we_nload_inst;
  wire plm_filters_rsc_req_vz_nload_inst;
  wire [66:0] dma_read_ctrl_rsc_dat_nload_inst;
  wire dma_read_ctrl_rsc_vld_nload_inst;
  wire dma_read_chnl_rsc_rdy_nload_inst;
  wire done_rsc_rdy_nload_inst;
  wire done_rsc_vld_nload_inst;
  wire plm_filters_rsc_we_nload_inst_buz;
  wire [255:0] conf_info_rsc_dat_ncompute_inst;
  wire conf_info_rsc_vld_ncompute_inst;
  wire conf_info_rsc_rdy_ncompute_inst;
  wire [13:0] plm_inputs_rsc_radr_ncompute_inst;
  wire [31:0] plm_inputs_rsc_q_ncompute_inst;
  wire plm_inputs_rsc_req_vz_ncompute_inst;
  wire [15:0] plm_filters_rsc_radr_ncompute_inst;
  wire [31:0] plm_filters_rsc_q_ncompute_inst;
  wire plm_filters_rsc_req_vz_ncompute_inst;
  wire [13:0] plm_outputs_rsc_wadr_ncompute_inst;
  wire [31:0] plm_outputs_rsc_d_ncompute_inst;
  wire plm_outputs_rsc_we_ncompute_inst;
  wire plm_outputs_rsc_req_vz_ncompute_inst;
  wire done_rsc_rdy_ncompute_inst;
  wire done_rsc_vld_ncompute_inst;
  wire plm_outputs_rsc_we_ncompute_inst_buz;
  wire [255:0] conf_info_rsc_dat_nstore_inst;
  wire conf_info_rsc_vld_nstore_inst;
  wire conf_info_rsc_rdy_nstore_inst;
  wire [13:0] plm_outputs_rsc_radr_nstore_inst;
  wire [31:0] plm_outputs_rsc_q_nstore_inst;
  wire plm_outputs_rsc_req_vz_nstore_inst;
  wire [66:0] dma_write_ctrl_rsc_dat_nstore_inst;
  wire dma_write_ctrl_rsc_vld_nstore_inst;
  wire [63:0] dma_write_chnl_rsc_dat_nstore_inst;
  wire dma_write_chnl_rsc_vld_nstore_inst;
  wire done_rsc_rdy_nstore_inst;
  wire done_rsc_vld_nstore_inst;
  wire config_done_cns_vld_nconv2d_cxx_catapult_core_inst;
  wire load_done_cns_vld_nconv2d_cxx_catapult_core_inst;
  wire compute_done_cns_vld_nconv2d_cxx_catapult_core_inst;
  wire store_done_cns_vld_nconv2d_cxx_catapult_core_inst;
  wire conf_info_rsc_rdy_nconfig_inst_bud;
  wire plm_conf_load_rsc_vld_nconfig_inst_bud;
  wire conf_info_rsc_rdy_nload_inst_bud;
  wire plm_conf_compute_rsc_vld_nconfig_inst_bud;
  wire conf_info_rsc_rdy_ncompute_inst_bud;
  wire plm_conf_store_rsc_vld_nconfig_inst_bud;
  wire conf_info_rsc_rdy_nstore_inst_bud;
  wire done_rsc_vld_nconfig_inst_bud;
  wire config_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud;
  wire plm_inputs_rsc_rls_lz_nload_inst_bud;
  wire plm_inputs_rsc_rls_lz_ncompute_inst_bud;
  wire plm_filters_rsc_we_nload_inst_buz_bud;
  wire plm_filters_rsc_rls_lz_nload_inst_bud;
  wire plm_filters_rsc_rls_lz_ncompute_inst_bud;
  wire dma_read_ctrl_rsc_vld_nload_inst_bud;
  wire dma_read_chnl_rsc_rdy_nload_inst_bud;
  wire done_rsc_vld_nload_inst_bud;
  wire load_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud;
  wire plm_outputs_rsc_we_ncompute_inst_buz_bud;
  wire plm_outputs_rsc_rls_lz_ncompute_inst_bud;
  wire plm_outputs_rsc_rls_lz_nstore_inst_bud;
  wire done_rsc_vld_ncompute_inst_bud;
  wire compute_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud;
  wire dma_write_ctrl_rsc_vld_nstore_inst_bud;
  wire dma_write_chnl_rsc_vld_nstore_inst_bud;
  wire done_rsc_vld_nstore_inst_bud;
  wire store_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud;
  wire acc_done_rsc_vld_nconv2d_cxx_catapult_core_inst_bud;
  wire plm_conf_load_unc_2;
  wire plm_conf_load_idle;
  wire plm_conf_compute_unc_2;
  wire plm_conf_compute_idle;
  wire plm_conf_store_unc_2;
  wire plm_conf_store_idle;
  wire plm_inputs_cns_R0;
  wire plm_inputs_cns_S1;
  wire plm_inputs_cns_R1;
  wire [31:0] plm_inputs_cns_d_shi0;
  wire [31:0] plm_inputs_cns_d_shi1;
  wire [31:0] plm_inputs_cns_q_sho0;
  wire [31:0] plm_inputs_cns_q_sho1;
  wire [13:0] plm_inputs_cns_radr_shi0;
  wire [13:0] plm_inputs_cns_radr_shi1;
  wire [13:0] plm_inputs_cns_wadr_shi0;
  wire [13:0] plm_inputs_cns_wadr_shi1;
  wire plm_inputs_cns_we_shi0;
  wire plm_inputs_cns_we_shi1;
  wire plm_filters_cns_R0;
  wire plm_filters_cns_S1;
  wire plm_filters_cns_R1;
  wire [31:0] plm_filters_cns_d_shi0;
  wire [31:0] plm_filters_cns_d_shi1;
  wire [31:0] plm_filters_cns_q_sho0;
  wire [31:0] plm_filters_cns_q_sho1;
  wire [15:0] plm_filters_cns_radr_shi0;
  wire [15:0] plm_filters_cns_radr_shi1;
  wire [15:0] plm_filters_cns_wadr_shi0;
  wire [15:0] plm_filters_cns_wadr_shi1;
  wire plm_filters_cns_we_shi0;
  wire plm_filters_cns_we_shi1;
  wire plm_outputs_cns_R0;
  wire plm_outputs_cns_S1;
  wire plm_outputs_cns_R1;
  wire [31:0] plm_outputs_cns_d_shi0;
  wire [31:0] plm_outputs_cns_d_shi1;
  wire [31:0] plm_outputs_cns_q_sho0;
  wire [31:0] plm_outputs_cns_q_sho1;
  wire [13:0] plm_outputs_cns_radr_shi0;
  wire [13:0] plm_outputs_cns_radr_shi1;
  wire [13:0] plm_outputs_cns_wadr_shi0;
  wire [13:0] plm_outputs_cns_wadr_shi1;
  wire plm_outputs_cns_we_shi0;
  wire plm_outputs_cns_we_shi1;
  wire plm_inputs_cns_S0_iff;
  wire plm_filters_rsc_we_nload_inst_buz_iff;
  wire plm_filters_rsc_we_nload_inst_buz_bud_iff;
  wire plm_filters_cns_S0_iff;
  wire plm_outputs_rsc_we_ncompute_inst_buz_iff;
  wire plm_outputs_rsc_we_ncompute_inst_buz_bud_iff;
  wire plm_outputs_cns_S0_iff;
  wire plm_inputs_cns_S0_dmo;
  wire plm_filters_cns_S0_dmo;
  wire plm_outputs_cns_S0_dmo;


  // Interconnect Declarations for Component Instantiations 
  wire [255:0] nl_config_inst_conf_info_rsc_dat;
  assign nl_config_inst_conf_info_rsc_dat = {conf_info_rsc_dat_batch , conf_info_rsc_dat_n_w
      , conf_info_rsc_dat_n_h , conf_info_rsc_dat_n_c , conf_info_rsc_dat_kern ,
      conf_info_rsc_dat_filt , conf_info_rsc_dat_same , conf_info_rsc_dat_stride};
  esp_acc_conv2d_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd38),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_conf_load_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_conf_load_rsc_rdy_nconfig_inst),
      .din_vld(plm_conf_load_rsc_vld_nconfig_inst_bud),
      .din(plm_conf_load_rsc_dat_nconfig_inst),
      .dout_rdy(conf_info_rsc_rdy_nload_inst),
      .dout_vld(conf_info_rsc_vld_nload_inst),
      .dout(conf_info_rsc_dat_nload_inst),
      .sz(plm_conf_load_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_conf_load_idle)
    );
  esp_acc_conv2d_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd39),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd4),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_conf_compute_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_conf_compute_rsc_rdy_nconfig_inst),
      .din_vld(plm_conf_compute_rsc_vld_nconfig_inst_bud),
      .din(plm_conf_compute_rsc_dat_nconfig_inst),
      .dout_rdy(conf_info_rsc_rdy_ncompute_inst),
      .dout_vld(conf_info_rsc_vld_ncompute_inst),
      .dout(conf_info_rsc_dat_ncompute_inst),
      .sz(plm_conf_compute_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_conf_compute_idle)
    );
  esp_acc_conv2d_cxx_catapult_ccs_pipe_v5 #(.rscid(32'sd40),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd4),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_conf_store_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_conf_store_rsc_rdy_nconfig_inst),
      .din_vld(plm_conf_store_rsc_vld_nconfig_inst_bud),
      .din(plm_conf_store_rsc_dat_nconfig_inst),
      .dout_rdy(conf_info_rsc_rdy_nstore_inst),
      .dout_vld(conf_info_rsc_vld_nstore_inst),
      .dout(conf_info_rsc_dat_nstore_inst),
      .sz(plm_conf_store_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_conf_store_idle)
    );
  esp_acc_conv2d_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd41)) config_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_nconfig_inst_bud),
      .dout_vld(done_rsc_rdy_nconfig_inst),
      .din_vld(config_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .din_rdy(config_done_cns_vld_nconv2d_cxx_catapult_core_inst)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd14),
  .data_width(32'sd32),
  .depth(32'sd10368),
  .latency(32'sd1)) plm_inputs_cns_comp (
      .clk(clk),
      .clken(1'b1),
      .d(plm_inputs_cns_d_shi0),
      .q(plm_inputs_cns_q_sho0),
      .radr(plm_inputs_cns_radr_shi0),
      .wadr(plm_inputs_cns_wadr_shi0),
      .we(plm_inputs_cns_we_shi0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd14),
  .data_width(32'sd32),
  .depth(32'sd10368),
  .latency(32'sd1)) plm_inputs_cns_comp_1 (
      .clk(clk),
      .clken(1'b1),
      .d(plm_inputs_cns_d_shi1),
      .q(plm_inputs_cns_q_sho1),
      .radr(plm_inputs_cns_radr_shi1),
      .wadr(plm_inputs_cns_wadr_shi1),
      .we(plm_inputs_cns_we_shi1)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd16),
  .data_width(32'sd32),
  .depth(32'sd50176),
  .latency(32'sd1)) plm_filters_cns_comp (
      .clk(clk),
      .clken(1'b1),
      .d(plm_filters_cns_d_shi0),
      .q(plm_filters_cns_q_sho0),
      .radr(plm_filters_cns_radr_shi0),
      .wadr(plm_filters_cns_wadr_shi0),
      .we(plm_filters_cns_we_shi0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd16),
  .data_width(32'sd32),
  .depth(32'sd50176),
  .latency(32'sd1)) plm_filters_cns_comp_1 (
      .clk(clk),
      .clken(1'b1),
      .d(plm_filters_cns_d_shi1),
      .q(plm_filters_cns_q_sho1),
      .radr(plm_filters_cns_radr_shi1),
      .wadr(plm_filters_cns_wadr_shi1),
      .we(plm_filters_cns_we_shi1)
    );
  esp_acc_conv2d_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd42)) load_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_nload_inst),
      .dout_vld(done_rsc_rdy_nload_inst),
      .din_vld(load_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .din_rdy(load_done_cns_vld_nconv2d_cxx_catapult_core_inst)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd14),
  .data_width(32'sd32),
  .depth(32'sd10368),
  .latency(32'sd1)) plm_outputs_cns_comp (
      .clk(clk),
      .clken(1'b1),
      .d(plm_outputs_cns_d_shi0),
      .q(plm_outputs_cns_q_sho0),
      .radr(plm_outputs_cns_radr_shi0),
      .wadr(plm_outputs_cns_wadr_shi0),
      .we(plm_outputs_cns_we_shi0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd14),
  .data_width(32'sd32),
  .depth(32'sd10368),
  .latency(32'sd1)) plm_outputs_cns_comp_1 (
      .clk(clk),
      .clken(1'b1),
      .d(plm_outputs_cns_d_shi1),
      .q(plm_outputs_cns_q_sho1),
      .radr(plm_outputs_cns_radr_shi1),
      .wadr(plm_outputs_cns_wadr_shi1),
      .we(plm_outputs_cns_we_shi1)
    );
  esp_acc_conv2d_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd43)) compute_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_ncompute_inst),
      .dout_vld(done_rsc_rdy_ncompute_inst),
      .din_vld(compute_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .din_rdy(compute_done_cns_vld_nconv2d_cxx_catapult_core_inst)
    );
  esp_acc_conv2d_cxx_catapult_ccs_sync_pipe_v1 #(.rscid(32'sd44)) store_done_cns_pipe
      (
      .dout_rdy(done_rsc_vld_nstore_inst),
      .dout_vld(done_rsc_rdy_nstore_inst),
      .din_vld(store_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .din_rdy(store_done_cns_vld_nconv2d_cxx_catapult_core_inst)
    );
  esp_acc_conv2d_cxx_catapult_config config_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(nl_config_inst_conf_info_rsc_dat[255:0]),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_nconfig_inst_bud),
      .plm_conf_load_rsc_dat(plm_conf_load_rsc_dat_nconfig_inst),
      .plm_conf_load_rsc_vld(plm_conf_load_rsc_vld_nconfig_inst_bud),
      .plm_conf_load_rsc_rdy(plm_conf_load_rsc_rdy_nconfig_inst),
      .plm_conf_compute_rsc_dat(plm_conf_compute_rsc_dat_nconfig_inst),
      .plm_conf_compute_rsc_vld(plm_conf_compute_rsc_vld_nconfig_inst_bud),
      .plm_conf_compute_rsc_rdy(plm_conf_compute_rsc_rdy_nconfig_inst),
      .plm_conf_store_rsc_dat(plm_conf_store_rsc_dat_nconfig_inst),
      .plm_conf_store_rsc_vld(plm_conf_store_rsc_vld_nconfig_inst_bud),
      .plm_conf_store_rsc_rdy(plm_conf_store_rsc_rdy_nconfig_inst),
      .done_rsc_rdy(done_rsc_rdy_nconfig_inst),
      .done_rsc_vld(done_rsc_vld_nconfig_inst_bud)
    );
  esp_acc_conv2d_cxx_catapult_load load_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat_nload_inst),
      .conf_info_rsc_vld(conf_info_rsc_vld_nload_inst),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_nload_inst_bud),
      .plm_inputs_rsc_wadr(plm_inputs_rsc_wadr_nload_inst),
      .plm_inputs_rsc_d(plm_inputs_rsc_d_nload_inst),
      .plm_inputs_rsc_we(plm_inputs_rsc_we_nload_inst),
      .plm_inputs_rsc_req_vz(plm_inputs_rsc_req_vz_nload_inst),
      .plm_inputs_rsc_rls_lz(plm_inputs_rsc_rls_lz_nload_inst_bud),
      .plm_filters_rsc_wadr(plm_filters_rsc_wadr_nload_inst),
      .plm_filters_rsc_d(plm_filters_rsc_d_nload_inst),
      .plm_filters_rsc_we(plm_filters_rsc_we_nload_inst),
      .plm_filters_rsc_req_vz(plm_filters_rsc_req_vz_nload_inst),
      .plm_filters_rsc_rls_lz(plm_filters_rsc_rls_lz_nload_inst_bud),
      .dma_read_ctrl_rsc_dat(dma_read_ctrl_rsc_dat_nload_inst),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld_nload_inst_bud),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy_nload_inst_bud),
      .done_rsc_rdy(done_rsc_rdy_nload_inst),
      .done_rsc_vld(done_rsc_vld_nload_inst_bud)
    );
  esp_acc_conv2d_cxx_catapult_compute compute_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat_ncompute_inst),
      .conf_info_rsc_vld(conf_info_rsc_vld_ncompute_inst),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_ncompute_inst_bud),
      .plm_inputs_rsc_radr(plm_inputs_rsc_radr_ncompute_inst),
      .plm_inputs_rsc_q(plm_inputs_rsc_q_ncompute_inst),
      .plm_inputs_rsc_req_vz(plm_inputs_rsc_req_vz_ncompute_inst),
      .plm_inputs_rsc_rls_lz(plm_inputs_rsc_rls_lz_ncompute_inst_bud),
      .plm_filters_rsc_radr(plm_filters_rsc_radr_ncompute_inst),
      .plm_filters_rsc_q(plm_filters_rsc_q_ncompute_inst),
      .plm_filters_rsc_req_vz(plm_filters_rsc_req_vz_ncompute_inst),
      .plm_filters_rsc_rls_lz(plm_filters_rsc_rls_lz_ncompute_inst_bud),
      .plm_outputs_rsc_wadr(plm_outputs_rsc_wadr_ncompute_inst),
      .plm_outputs_rsc_d(plm_outputs_rsc_d_ncompute_inst),
      .plm_outputs_rsc_we(plm_outputs_rsc_we_ncompute_inst),
      .plm_outputs_rsc_req_vz(plm_outputs_rsc_req_vz_ncompute_inst),
      .plm_outputs_rsc_rls_lz(plm_outputs_rsc_rls_lz_ncompute_inst_bud),
      .done_rsc_rdy(done_rsc_rdy_ncompute_inst),
      .done_rsc_vld(done_rsc_vld_ncompute_inst_bud)
    );
  esp_acc_conv2d_cxx_catapult_store store_inst (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat(conf_info_rsc_dat_nstore_inst),
      .conf_info_rsc_vld(conf_info_rsc_vld_nstore_inst),
      .conf_info_rsc_rdy(conf_info_rsc_rdy_nstore_inst_bud),
      .plm_outputs_rsc_radr(plm_outputs_rsc_radr_nstore_inst),
      .plm_outputs_rsc_q(plm_outputs_rsc_q_nstore_inst),
      .plm_outputs_rsc_req_vz(plm_outputs_rsc_req_vz_nstore_inst),
      .plm_outputs_rsc_rls_lz(plm_outputs_rsc_rls_lz_nstore_inst_bud),
      .dma_write_ctrl_rsc_dat(dma_write_ctrl_rsc_dat_nstore_inst),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld_nstore_inst_bud),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat_nstore_inst),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld_nstore_inst_bud),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .done_rsc_rdy(done_rsc_rdy_nstore_inst),
      .done_rsc_vld(done_rsc_vld_nstore_inst_bud)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_core conv2d_cxx_catapult_core_inst
      (
      .clk(clk),
      .rst(rst),
      .acc_done_rsc_vld(acc_done_rsc_vld_nconv2d_cxx_catapult_core_inst_bud),
      .config_done_cns_rdy(config_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .config_done_cns_vld(config_done_cns_vld_nconv2d_cxx_catapult_core_inst),
      .load_done_cns_rdy(load_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .load_done_cns_vld(load_done_cns_vld_nconv2d_cxx_catapult_core_inst),
      .compute_done_cns_rdy(compute_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .compute_done_cns_vld(compute_done_cns_vld_nconv2d_cxx_catapult_core_inst),
      .store_done_cns_rdy(store_done_cns_rdy_nconv2d_cxx_catapult_core_inst_bud),
      .store_done_cns_vld(store_done_cns_vld_nconv2d_cxx_catapult_core_inst)
    );
  esp_acc_conv2d_cxx_catapult_unreg_hier unreg (
      .in_0(plm_inputs_cns_S0_iff),
      .out_0(plm_inputs_cns_R0)
    );
  esp_acc_conv2d_cxx_catapult_unreg_hier unreg_1 (
      .in_0(plm_inputs_cns_S1),
      .out_0(plm_inputs_cns_R1)
    );
  esp_acc_conv2d_cxx_catapult_unreg_hier unreg_2 (
      .in_0(plm_filters_cns_S0_iff),
      .out_0(plm_filters_cns_R0)
    );
  esp_acc_conv2d_cxx_catapult_unreg_hier unreg_3 (
      .in_0(plm_filters_cns_S1),
      .out_0(plm_filters_cns_R1)
    );
  esp_acc_conv2d_cxx_catapult_unreg_hier unreg_4 (
      .in_0(plm_outputs_cns_S0_iff),
      .out_0(plm_outputs_cns_R0)
    );
  esp_acc_conv2d_cxx_catapult_unreg_hier unreg_5 (
      .in_0(plm_outputs_cns_S1),
      .out_0(plm_outputs_cns_R1)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_cKlrPsts_cns_bctl conv2d_cxx_cKlrPsts_cns_bctl_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_rdy_nload_inst(conf_info_rsc_rdy_nload_inst),
      .plm_inputs_rsc_wadr_nload_inst(plm_inputs_rsc_wadr_nload_inst),
      .plm_inputs_rsc_d_nload_inst(plm_inputs_rsc_d_nload_inst),
      .plm_inputs_rsc_we_nload_inst(plm_inputs_rsc_we_nload_inst),
      .plm_inputs_rsc_req_vz_nload_inst(plm_inputs_rsc_req_vz_nload_inst),
      .dma_read_ctrl_rsc_vld_nload_inst(dma_read_ctrl_rsc_vld_nload_inst),
      .dma_read_chnl_rsc_rdy_nload_inst(dma_read_chnl_rsc_rdy_nload_inst),
      .done_rsc_vld_nload_inst(done_rsc_vld_nload_inst),
      .plm_filters_rsc_we_nload_inst_buz(plm_filters_rsc_we_nload_inst_buz),
      .conf_info_rsc_rdy_ncompute_inst(conf_info_rsc_rdy_ncompute_inst),
      .plm_inputs_rsc_radr_ncompute_inst(plm_inputs_rsc_radr_ncompute_inst),
      .plm_inputs_rsc_q_ncompute_inst(plm_inputs_rsc_q_ncompute_inst),
      .plm_inputs_rsc_req_vz_ncompute_inst(plm_inputs_rsc_req_vz_ncompute_inst),
      .done_rsc_vld_ncompute_inst(done_rsc_vld_ncompute_inst),
      .plm_outputs_rsc_we_ncompute_inst_buz(plm_outputs_rsc_we_ncompute_inst_buz),
      .conf_info_rsc_rdy_nload_inst_bud(conf_info_rsc_rdy_nload_inst_bud),
      .conf_info_rsc_rdy_ncompute_inst_bud(conf_info_rsc_rdy_ncompute_inst_bud),
      .plm_inputs_rsc_rls_lz_nload_inst_bud(plm_inputs_rsc_rls_lz_nload_inst_bud),
      .plm_inputs_rsc_rls_lz_ncompute_inst_bud(plm_inputs_rsc_rls_lz_ncompute_inst_bud),
      .plm_filters_rsc_we_nload_inst_buz_bud(plm_filters_rsc_we_nload_inst_buz_bud),
      .plm_filters_rsc_rls_lz_nload_inst_bud(1'b0),
      .plm_filters_rsc_rls_lz_ncompute_inst_bud(1'b0),
      .dma_read_ctrl_rsc_vld_nload_inst_bud(dma_read_ctrl_rsc_vld_nload_inst_bud),
      .dma_read_chnl_rsc_rdy_nload_inst_bud(dma_read_chnl_rsc_rdy_nload_inst_bud),
      .done_rsc_vld_nload_inst_bud(done_rsc_vld_nload_inst_bud),
      .plm_outputs_rsc_we_ncompute_inst_buz_bud(plm_outputs_rsc_we_ncompute_inst_buz_bud),
      .plm_outputs_rsc_rls_lz_ncompute_inst_bud(1'b0),
      .done_rsc_vld_ncompute_inst_bud(done_rsc_vld_ncompute_inst_bud),
      .plm_inputs_cns_S0(plm_inputs_cns_S0_dmo),
      .plm_inputs_cns_R0(plm_inputs_cns_R0),
      .plm_inputs_cns_S1(plm_inputs_cns_S1),
      .plm_inputs_cns_R1(plm_inputs_cns_R1),
      .plm_inputs_cns_d_shi0(plm_inputs_cns_d_shi0),
      .plm_inputs_cns_d_shi1(plm_inputs_cns_d_shi1),
      .plm_inputs_cns_q_sho0(plm_inputs_cns_q_sho0),
      .plm_inputs_cns_q_sho1(plm_inputs_cns_q_sho1),
      .plm_inputs_cns_radr_shi0(plm_inputs_cns_radr_shi0),
      .plm_inputs_cns_radr_shi1(plm_inputs_cns_radr_shi1),
      .plm_inputs_cns_wadr_shi0(plm_inputs_cns_wadr_shi0),
      .plm_inputs_cns_wadr_shi1(plm_inputs_cns_wadr_shi1),
      .plm_inputs_cns_we_shi0(plm_inputs_cns_we_shi0),
      .plm_inputs_cns_we_shi1(plm_inputs_cns_we_shi1),
      .plm_inputs_cns_S0_pff(plm_inputs_cns_S0_iff),
      .plm_filters_rsc_we_nload_inst_buz_pff(plm_filters_rsc_we_nload_inst_buz_iff),
      .plm_filters_rsc_we_nload_inst_buz_bud_pff(plm_filters_rsc_we_nload_inst_buz_bud_iff),
      .plm_outputs_rsc_we_ncompute_inst_buz_pff(plm_outputs_rsc_we_ncompute_inst_buz_iff),
      .plm_outputs_rsc_we_ncompute_inst_buz_bud_pff(plm_outputs_rsc_we_ncompute_inst_buz_bud_iff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_cYDPQCrs_cns_bctl conv2d_cxx_cYDPQCrs_cns_bctl_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_filters_rsc_wadr_nload_inst(plm_filters_rsc_wadr_nload_inst),
      .plm_filters_rsc_d_nload_inst(plm_filters_rsc_d_nload_inst),
      .plm_filters_rsc_we_nload_inst(plm_filters_rsc_we_nload_inst),
      .plm_filters_rsc_req_vz_nload_inst(plm_filters_rsc_req_vz_nload_inst),
      .plm_filters_rsc_we_nload_inst_buz(1'b0),
      .plm_filters_rsc_radr_ncompute_inst(plm_filters_rsc_radr_ncompute_inst),
      .plm_filters_rsc_q_ncompute_inst(plm_filters_rsc_q_ncompute_inst),
      .plm_filters_rsc_req_vz_ncompute_inst(plm_filters_rsc_req_vz_ncompute_inst),
      .plm_filters_rsc_we_nload_inst_buz_bud(plm_filters_rsc_we_nload_inst_buz_bud),
      .plm_filters_rsc_rls_lz_nload_inst_bud(plm_filters_rsc_rls_lz_nload_inst_bud),
      .plm_filters_rsc_rls_lz_ncompute_inst_bud(plm_filters_rsc_rls_lz_ncompute_inst_bud),
      .plm_filters_cns_S0(plm_filters_cns_S0_dmo),
      .plm_filters_cns_R0(plm_filters_cns_R0),
      .plm_filters_cns_S1(plm_filters_cns_S1),
      .plm_filters_cns_R1(plm_filters_cns_R1),
      .plm_filters_cns_d_shi0(plm_filters_cns_d_shi0),
      .plm_filters_cns_d_shi1(plm_filters_cns_d_shi1),
      .plm_filters_cns_q_sho0(plm_filters_cns_q_sho0),
      .plm_filters_cns_q_sho1(plm_filters_cns_q_sho1),
      .plm_filters_cns_radr_shi0(plm_filters_cns_radr_shi0),
      .plm_filters_cns_radr_shi1(plm_filters_cns_radr_shi1),
      .plm_filters_cns_wadr_shi0(plm_filters_cns_wadr_shi0),
      .plm_filters_cns_wadr_shi1(plm_filters_cns_wadr_shi1),
      .plm_filters_cns_we_shi0(plm_filters_cns_we_shi0),
      .plm_filters_cns_we_shi1(plm_filters_cns_we_shi1),
      .plm_filters_rsc_we_nload_inst_buz_pff(plm_filters_rsc_we_nload_inst_buz_iff),
      .plm_filters_rsc_we_nload_inst_buz_bud_pff(plm_filters_rsc_we_nload_inst_buz_bud_iff),
      .plm_filters_cns_S0_pff(plm_filters_cns_S0_iff)
    );
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_cYqiuTts_cns_bctl conv2d_cxx_cYqiuTts_cns_bctl_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_outputs_rsc_wadr_ncompute_inst(plm_outputs_rsc_wadr_ncompute_inst),
      .plm_outputs_rsc_d_ncompute_inst(plm_outputs_rsc_d_ncompute_inst),
      .plm_outputs_rsc_we_ncompute_inst(plm_outputs_rsc_we_ncompute_inst),
      .plm_outputs_rsc_req_vz_ncompute_inst(plm_outputs_rsc_req_vz_ncompute_inst),
      .plm_outputs_rsc_we_ncompute_inst_buz(1'b0),
      .conf_info_rsc_rdy_nstore_inst(conf_info_rsc_rdy_nstore_inst),
      .plm_outputs_rsc_radr_nstore_inst(plm_outputs_rsc_radr_nstore_inst),
      .plm_outputs_rsc_q_nstore_inst(plm_outputs_rsc_q_nstore_inst),
      .plm_outputs_rsc_req_vz_nstore_inst(plm_outputs_rsc_req_vz_nstore_inst),
      .dma_write_ctrl_rsc_vld_nstore_inst(dma_write_ctrl_rsc_vld_nstore_inst),
      .dma_write_chnl_rsc_vld_nstore_inst(dma_write_chnl_rsc_vld_nstore_inst),
      .done_rsc_vld_nstore_inst(done_rsc_vld_nstore_inst),
      .conf_info_rsc_rdy_nstore_inst_bud(conf_info_rsc_rdy_nstore_inst_bud),
      .plm_outputs_rsc_we_ncompute_inst_buz_bud(plm_outputs_rsc_we_ncompute_inst_buz_bud),
      .plm_outputs_rsc_rls_lz_ncompute_inst_bud(plm_outputs_rsc_rls_lz_ncompute_inst_bud),
      .plm_outputs_rsc_rls_lz_nstore_inst_bud(plm_outputs_rsc_rls_lz_nstore_inst_bud),
      .dma_write_ctrl_rsc_vld_nstore_inst_bud(dma_write_ctrl_rsc_vld_nstore_inst_bud),
      .dma_write_chnl_rsc_vld_nstore_inst_bud(dma_write_chnl_rsc_vld_nstore_inst_bud),
      .done_rsc_vld_nstore_inst_bud(done_rsc_vld_nstore_inst_bud),
      .plm_outputs_cns_S0(plm_outputs_cns_S0_dmo),
      .plm_outputs_cns_R0(plm_outputs_cns_R0),
      .plm_outputs_cns_S1(plm_outputs_cns_S1),
      .plm_outputs_cns_R1(plm_outputs_cns_R1),
      .plm_outputs_cns_d_shi0(plm_outputs_cns_d_shi0),
      .plm_outputs_cns_d_shi1(plm_outputs_cns_d_shi1),
      .plm_outputs_cns_q_sho0(plm_outputs_cns_q_sho0),
      .plm_outputs_cns_q_sho1(plm_outputs_cns_q_sho1),
      .plm_outputs_cns_radr_shi0(plm_outputs_cns_radr_shi0),
      .plm_outputs_cns_radr_shi1(plm_outputs_cns_radr_shi1),
      .plm_outputs_cns_wadr_shi0(plm_outputs_cns_wadr_shi0),
      .plm_outputs_cns_wadr_shi1(plm_outputs_cns_wadr_shi1),
      .plm_outputs_cns_we_shi0(plm_outputs_cns_we_shi0),
      .plm_outputs_cns_we_shi1(plm_outputs_cns_we_shi1),
      .plm_outputs_rsc_we_ncompute_inst_buz_pff(plm_outputs_rsc_we_ncompute_inst_buz_iff),
      .plm_outputs_rsc_we_ncompute_inst_buz_bud_pff(plm_outputs_rsc_we_ncompute_inst_buz_bud_iff),
      .plm_outputs_cns_S0_pff(plm_outputs_cns_S0_iff)
    );
  assign conf_info_rsc_rdy = conf_info_rsc_rdy_nconfig_inst_bud;
  assign dma_read_ctrl_rsc_dat_index = dma_read_ctrl_rsc_dat_nload_inst[31:0];
  assign dma_read_ctrl_rsc_dat_length = dma_read_ctrl_rsc_dat_nload_inst[63:32];
  assign dma_read_ctrl_rsc_dat_size = dma_read_ctrl_rsc_dat_nload_inst[66:64];
  assign dma_write_ctrl_rsc_dat_index = dma_write_ctrl_rsc_dat_nstore_inst[31:0];
  assign dma_write_ctrl_rsc_dat_length = dma_write_ctrl_rsc_dat_nstore_inst[63:32];
  assign dma_write_ctrl_rsc_dat_size = dma_write_ctrl_rsc_dat_nstore_inst[66:64];
  assign dma_read_ctrl_rsc_vld = dma_read_ctrl_rsc_vld_nload_inst;
  assign dma_read_chnl_rsc_rdy = dma_read_chnl_rsc_rdy_nload_inst;
  assign dma_write_ctrl_rsc_vld = dma_write_ctrl_rsc_vld_nstore_inst;
  assign dma_write_chnl_rsc_vld = dma_write_chnl_rsc_vld_nstore_inst;
  assign dma_write_chnl_rsc_dat = dma_write_chnl_rsc_dat_nstore_inst;
  assign acc_done_rsc_vld = acc_done_rsc_vld_nconv2d_cxx_catapult_core_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    conv2d_cxx_catapult_hier_fx32_dma64
// ------------------------------------------------------------------


module conv2d_cxx_catapult_hier_fx32_dma64 (
  clk, rst, conf_info_rsc_dat, conf_info_rsc_vld, conf_info_rsc_rdy, dma_read_ctrl_rsc_dat,
      dma_read_ctrl_rsc_vld, dma_read_ctrl_rsc_rdy, dma_write_ctrl_rsc_dat, dma_write_ctrl_rsc_vld,
      dma_write_ctrl_rsc_rdy, dma_read_chnl_rsc_dat, dma_read_chnl_rsc_vld, dma_read_chnl_rsc_rdy,
      dma_write_chnl_rsc_dat, dma_write_chnl_rsc_vld, dma_write_chnl_rsc_rdy, acc_done_rsc_vld
);
  input clk;
  input rst;
  input [255:0] conf_info_rsc_dat;
  input conf_info_rsc_vld;
  output conf_info_rsc_rdy;
  output [66:0] dma_read_ctrl_rsc_dat;
  output dma_read_ctrl_rsc_vld;
  input dma_read_ctrl_rsc_rdy;
  output [66:0] dma_write_ctrl_rsc_dat;
  output dma_write_ctrl_rsc_vld;
  input dma_write_ctrl_rsc_rdy;
  input [63:0] dma_read_chnl_rsc_dat;
  input dma_read_chnl_rsc_vld;
  output dma_read_chnl_rsc_rdy;
  output [63:0] dma_write_chnl_rsc_dat;
  output dma_write_chnl_rsc_vld;
  input dma_write_chnl_rsc_rdy;
  output acc_done_rsc_vld;


  // Interconnect Declarations
  wire [2:0] dma_read_ctrl_rsc_dat_size;
  wire [31:0] dma_read_ctrl_rsc_dat_length;
  wire [31:0] dma_read_ctrl_rsc_dat_index;
  wire [2:0] dma_write_ctrl_rsc_dat_size;
  wire [31:0] dma_write_ctrl_rsc_dat_length;
  wire [31:0] dma_write_ctrl_rsc_dat_index;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_batch;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_batch = conf_info_rsc_dat[255:224];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w = conf_info_rsc_dat[223:192];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h = conf_info_rsc_dat[191:160];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c = conf_info_rsc_dat[159:128];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_kern;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_kern = conf_info_rsc_dat[127:96];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_filt;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_filt = conf_info_rsc_dat[95:64];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_same;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_same = conf_info_rsc_dat[63:32];
  wire [31:0] nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_stride;
  assign nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_stride = conf_info_rsc_dat[31:0];
  esp_acc_conv2d_cxx_catapult_conv2d_cxx_catapult_struct conv2d_cxx_catapult_struct_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info_rsc_dat_batch(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_batch[31:0]),
      .conf_info_rsc_dat_n_w(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_w[31:0]),
      .conf_info_rsc_dat_n_h(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_h[31:0]),
      .conf_info_rsc_dat_n_c(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_n_c[31:0]),
      .conf_info_rsc_dat_kern(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_kern[31:0]),
      .conf_info_rsc_dat_filt(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_filt[31:0]),
      .conf_info_rsc_dat_same(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_same[31:0]),
      .conf_info_rsc_dat_stride(nl_conv2d_cxx_catapult_struct_inst_conf_info_rsc_dat_stride[31:0]),
      .conf_info_rsc_vld(conf_info_rsc_vld),
      .conf_info_rsc_rdy(conf_info_rsc_rdy),
      .dma_read_ctrl_rsc_dat_size(dma_read_ctrl_rsc_dat_size),
      .dma_read_ctrl_rsc_dat_length(dma_read_ctrl_rsc_dat_length),
      .dma_read_ctrl_rsc_dat_index(dma_read_ctrl_rsc_dat_index),
      .dma_read_ctrl_rsc_vld(dma_read_ctrl_rsc_vld),
      .dma_read_ctrl_rsc_rdy(dma_read_ctrl_rsc_rdy),
      .dma_write_ctrl_rsc_dat_size(dma_write_ctrl_rsc_dat_size),
      .dma_write_ctrl_rsc_dat_length(dma_write_ctrl_rsc_dat_length),
      .dma_write_ctrl_rsc_dat_index(dma_write_ctrl_rsc_dat_index),
      .dma_write_ctrl_rsc_vld(dma_write_ctrl_rsc_vld),
      .dma_write_ctrl_rsc_rdy(dma_write_ctrl_rsc_rdy),
      .dma_read_chnl_rsc_dat(dma_read_chnl_rsc_dat),
      .dma_read_chnl_rsc_vld(dma_read_chnl_rsc_vld),
      .dma_read_chnl_rsc_rdy(dma_read_chnl_rsc_rdy),
      .dma_write_chnl_rsc_dat(dma_write_chnl_rsc_dat),
      .dma_write_chnl_rsc_vld(dma_write_chnl_rsc_vld),
      .dma_write_chnl_rsc_rdy(dma_write_chnl_rsc_rdy),
      .acc_done_rsc_vld(acc_done_rsc_vld)
    );
  assign dma_read_ctrl_rsc_dat = {dma_read_ctrl_rsc_dat_size , dma_read_ctrl_rsc_dat_length
      , dma_read_ctrl_rsc_dat_index};
  assign dma_write_ctrl_rsc_dat = {dma_write_ctrl_rsc_dat_size , dma_write_ctrl_rsc_dat_length
      , dma_write_ctrl_rsc_dat_index};
endmodule



